.SUBCKT not1 A VDD VSS ZN 
M_M1 N_ZN_M0_d N_A_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.028350P PS=0.750000U PD=0.750000U
M_M0 N_ZN_M1_d N_A_M1_g N_VSS_M1_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.018900P PS=0.570000U PD=0.570000U
C_x_PM_INV_X2__VSS_c0 VSS VSS 4.27233e-17
C_x_PM_INV_X2__VSS_c1 VSS x_PM_INV_X2__VSS_6 1.03058e-17
C_x_PM_INV_X2__VSS_c2 VSS N_VSS_M1_s 1.41503e-17
R_x_PM_INV_X2__VSS_r3 VSS x_PM_INV_X2__VSS_6 0.178824
R_x_PM_INV_X2__VSS_r4 x_PM_INV_X2__VSS_6 x_PM_INV_X2__VSS_2 0.264221
R_x_PM_INV_X2__VSS_r5 N_VSS_M1_s x_PM_INV_X2__VSS_2 0.230714
C_x_PM_INV_X2__VDD_c0 VSS VDD 4.06353e-17
C_x_PM_INV_X2__VDD_c1 VSS N_VDD_M0_s 3.31015e-17
C_x_PM_INV_X2__VDD_c2 VSS x_PM_INV_X2__VDD_2 1.05089e-17
R_x_PM_INV_X2__VDD_r3 VDD x_PM_INV_X2__VDD_2 0.0689273
R_x_PM_INV_X2__VDD_r4 N_VDD_M0_s x_PM_INV_X2__VDD_2 0.420714
C_x_PM_INV_X2__A_c0 VSS x_PM_INV_X2__A_14 8.49814e-18
C_x_PM_INV_X2__A_c1 VSS x_PM_INV_X2__A_12 3.56395e-17
C_x_PM_INV_X2__A_c2 VSS N_A_M0_g 9.12771e-17
C_x_PM_INV_X2__A_c3 VSS N_A_M1_g 4.61923e-17
R_x_PM_INV_X2__A_r4 x_PM_INV_X2__A_18 x_PM_INV_X2__A_14 4.74714
R_x_PM_INV_X2__A_r5 x_PM_INV_X2__A_17 x_PM_INV_X2__A_14 4.74714
R_x_PM_INV_X2__A_r6 x_PM_INV_X2__A_14 x_PM_INV_X2__A_12 25.0012
R_x_PM_INV_X2__A_r7 x_PM_INV_X2__A_12 A 0.156071
R_x_PM_INV_X2__A_r8 N_A_M0_g x_PM_INV_X2__A_18 95.94
R_x_PM_INV_X2__A_r9 N_A_M1_g x_PM_INV_X2__A_17 42.12
C_x_PM_INV_X2__ZN_c0 VSS N_ZN_M1_d 3.90212e-17
C_x_PM_INV_X2__ZN_c1 VSS ZN 7.52075e-17
C_x_PM_INV_X2__ZN_c2 VSS N_ZN_M0_d 5.26306e-17
C_x_PM_INV_X2__ZN_c3 VSS x_PM_INV_X2__ZN_3 4.60415e-18
R_x_PM_INV_X2__ZN_r4 ZN x_PM_INV_X2__ZN_8 1.87286
R_x_PM_INV_X2__ZN_r5 x_PM_INV_X2__ZN_7 N_ZN_M1_d 0.30478
R_x_PM_INV_X2__ZN_r6 ZN x_PM_INV_X2__ZN_7 1.87286
R_x_PM_INV_X2__ZN_r7 x_PM_INV_X2__ZN_8 x_PM_INV_X2__ZN_3 0.20978
R_x_PM_INV_X2__ZN_r8 N_ZN_M0_d x_PM_INV_X2__ZN_3 0.686111
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
