
module c880_tb();

reg N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

wire N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

	 
c880 c0(N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
		 N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
		 N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
		 N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
		 N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
		 N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
		 N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
		 N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
		 N865,N866,N874,N878,N879,N880);
		 
	 
reg [59:0] test_vectors[0:9];	
reg [25:0] out_vectors[0:9];	

integer k;
			 
initial
	begin

	$readmemb("c880_input_data.txt", test_vectors);
	
	end
	
initial
	begin
	
	for(k = 0; k < 10; k = k + 1)
		begin		
		#10
		{N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268} = test_vectors[k];
			
		#1
		out_vectors[k] = {N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880};
		 
		$display("output%d: %h\n", k, out_vectors[k]);
		
		end
		
		$writememb("c880_in_data.txt", test_vectors);
		$writememb("c880_out_data.txt", out_vectors);
	
	end



endmodule
