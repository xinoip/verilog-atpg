.SUBCKT nor4 A1 A2 A3 A4 VDD VSS ZN
M_M4 8 N_A4_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.650000U AS=0.068250P AD=0.091000P PS=1.510000U PD=1.580000U
M_M5 9 N_A3_M1_g 8 VDD PMOS_VTL L=0.050U W=0.650000U AS=0.091000P AD=0.091000P PS=1.580000U PD=1.580000U
M_M6 10 N_A2_M2_g 9 VDD PMOS_VTL L=0.050U W=0.650000U AS=0.091000P AD=0.091000P PS=1.580000U PD=1.580000U
M_M7 N_ZN_M3_d N_A1_M3_g 10 VDD PMOS_VTL L=0.050U W=0.650000U AS=0.091000P AD=0.068250P PS=1.580000U PD=1.510000U
M_M0 N_ZN_M4_d N_A4_M4_g N_VSS_M4_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M_M1 N_VSS_M5_d N_A3_M5_g N_ZN_M4_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M_M2 N_ZN_M6_d N_A2_M6_g N_VSS_M5_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M_M3 N_VSS_M7_d N_A1_M7_g N_ZN_M6_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_NOR4_X2__VSS_c0 VSS VSS 2.64443e-18
C_x_PM_NOR4_X2__VSS_c1 VSS N_VSS_M7_d 1.30717e-17
C_x_PM_NOR4_X2__VSS_c2 VSS x_PM_NOR4_X2__VSS_14 5.3438e-17
C_x_PM_NOR4_X2__VSS_c3 VSS N_VSS_M5_d 2.04204e-17
C_x_PM_NOR4_X2__VSS_c4 VSS x_PM_NOR4_X2__VSS_9 1.06295e-17
C_x_PM_NOR4_X2__VSS_c5 VSS x_PM_NOR4_X2__VSS_8 3.88904e-17
C_x_PM_NOR4_X2__VSS_c6 VSS N_VSS_M4_s 1.0831e-17
R_x_PM_NOR4_X2__VSS_r7 N_VSS_M7_d x_PM_NOR4_X2__VSS_16 0.230714
R_x_PM_NOR4_X2__VSS_r8 VSS x_PM_NOR4_X2__VSS_15 0.0731438
R_x_PM_NOR4_X2__VSS_r9 x_PM_NOR4_X2__VSS_16 x_PM_NOR4_X2__VSS_14 0.264221
R_x_PM_NOR4_X2__VSS_r10 x_PM_NOR4_X2__VSS_15 x_PM_NOR4_X2__VSS_14 0.681765
R_x_PM_NOR4_X2__VSS_r11 VSS x_PM_NOR4_X2__VSS_10 0.145286
R_x_PM_NOR4_X2__VSS_r12 N_VSS_M5_d x_PM_NOR4_X2__VSS_10 0.230714
R_x_PM_NOR4_X2__VSS_r13 VSS x_PM_NOR4_X2__VSS_8 0.0731438
R_x_PM_NOR4_X2__VSS_r14 x_PM_NOR4_X2__VSS_9 x_PM_NOR4_X2__VSS_8 0.692941
R_x_PM_NOR4_X2__VSS_r15 x_PM_NOR4_X2__VSS_9 x_PM_NOR4_X2__VSS_4 0.264221
R_x_PM_NOR4_X2__VSS_r16 N_VSS_M4_s x_PM_NOR4_X2__VSS_4 0.230714
C_x_PM_NOR4_X2__VDD_c0 VSS VDD 7.40695e-17
C_x_PM_NOR4_X2__VDD_c1 VSS N_VDD_M0_s 2.4691e-17
C_x_PM_NOR4_X2__VDD_c2 VSS x_PM_NOR4_X2__VDD_2 1.06862e-17
R_x_PM_NOR4_X2__VDD_r3 VDD x_PM_NOR4_X2__VDD_2 0.0689273
R_x_PM_NOR4_X2__VDD_r4 N_VDD_M0_s x_PM_NOR4_X2__VDD_2 0.230714
C_x_PM_NOR4_X2__A4_c0 VSS x_PM_NOR4_X2__A4_14 7.18659e-18
C_x_PM_NOR4_X2__A4_c1 VSS x_PM_NOR4_X2__A4_12 3.56769e-17
C_x_PM_NOR4_X2__A4_c2 VSS N_A4_M0_g 7.98018e-17
C_x_PM_NOR4_X2__A4_c3 VSS N_A4_M4_g 4.23053e-17
R_x_PM_NOR4_X2__A4_r4 x_PM_NOR4_X2__A4_18 x_PM_NOR4_X2__A4_14 4.74714
R_x_PM_NOR4_X2__A4_r5 x_PM_NOR4_X2__A4_17 x_PM_NOR4_X2__A4_14 4.74714
R_x_PM_NOR4_X2__A4_r6 x_PM_NOR4_X2__A4_14 x_PM_NOR4_X2__A4_12 25.0012
R_x_PM_NOR4_X2__A4_r7 x_PM_NOR4_X2__A4_12 A4 0.156071
R_x_PM_NOR4_X2__A4_r8 N_A4_M0_g x_PM_NOR4_X2__A4_18 70.98
R_x_PM_NOR4_X2__A4_r9 N_A4_M4_g x_PM_NOR4_X2__A4_17 42.9
C_x_PM_NOR4_X2__ZN_c0 VSS x_PM_NOR4_X2__ZN_27 1.32309e-17
C_x_PM_NOR4_X2__ZN_c1 VSS x_PM_NOR4_X2__ZN_26 2.32902e-17
C_x_PM_NOR4_X2__ZN_c2 VSS x_PM_NOR4_X2__ZN_23 4.60612e-17
C_x_PM_NOR4_X2__ZN_c3 VSS N_ZN_M3_d 2.50235e-17
C_x_PM_NOR4_X2__ZN_c4 VSS x_PM_NOR4_X2__ZN_18 3.46798e-18
C_x_PM_NOR4_X2__ZN_c5 VSS x_PM_NOR4_X2__ZN_16 2.65091e-17
C_x_PM_NOR4_X2__ZN_c6 VSS N_ZN_M6_d 2.42211e-17
C_x_PM_NOR4_X2__ZN_c7 VSS x_PM_NOR4_X2__ZN_11 2.27649e-17
C_x_PM_NOR4_X2__ZN_c8 VSS x_PM_NOR4_X2__ZN_10 1.9661e-17
C_x_PM_NOR4_X2__ZN_c9 VSS x_PM_NOR4_X2__ZN_9 1.62159e-17
C_x_PM_NOR4_X2__ZN_c10 VSS N_ZN_M4_d 2.33665e-17
R_x_PM_NOR4_X2__ZN_r11 x_PM_NOR4_X2__ZN_26 ZN 0.189936
R_x_PM_NOR4_X2__ZN_r12 x_PM_NOR4_X2__ZN_23 x_PM_NOR4_X2__ZN_22 1.65571
R_x_PM_NOR4_X2__ZN_r13 x_PM_NOR4_X2__ZN_23 x_PM_NOR4_X2__ZN_18 0.192227
R_x_PM_NOR4_X2__ZN_r14 N_ZN_M3_d x_PM_NOR4_X2__ZN_18 0.861333
R_x_PM_NOR4_X2__ZN_r15 x_PM_NOR4_X2__ZN_27 x_PM_NOR4_X2__ZN_17 0.113465
R_x_PM_NOR4_X2__ZN_r16 x_PM_NOR4_X2__ZN_22 x_PM_NOR4_X2__ZN_16 0.212317
R_x_PM_NOR4_X2__ZN_r17 x_PM_NOR4_X2__ZN_17 x_PM_NOR4_X2__ZN_16 0.705714
R_x_PM_NOR4_X2__ZN_r18 x_PM_NOR4_X2__ZN_27 x_PM_NOR4_X2__ZN_12 0.0883294
R_x_PM_NOR4_X2__ZN_r19 N_ZN_M6_d x_PM_NOR4_X2__ZN_12 0.257857
R_x_PM_NOR4_X2__ZN_r20 ZN x_PM_NOR4_X2__ZN_11 0.095
R_x_PM_NOR4_X2__ZN_r21 x_PM_NOR4_X2__ZN_27 x_PM_NOR4_X2__ZN_10 0.113465
R_x_PM_NOR4_X2__ZN_r22 x_PM_NOR4_X2__ZN_11 x_PM_NOR4_X2__ZN_10 0.257857
R_x_PM_NOR4_X2__ZN_r23 x_PM_NOR4_X2__ZN_9 x_PM_NOR4_X2__ZN_26 0.732857
R_x_PM_NOR4_X2__ZN_r24 x_PM_NOR4_X2__ZN_9 x_PM_NOR4_X2__ZN_4 0.212317
R_x_PM_NOR4_X2__ZN_r25 N_ZN_M4_d x_PM_NOR4_X2__ZN_4 0.257857
C_x_PM_NOR4_X2__A3_c0 VSS x_PM_NOR4_X2__A3_14 8.988e-18
C_x_PM_NOR4_X2__A3_c1 VSS x_PM_NOR4_X2__A3_12 6.21612e-17
C_x_PM_NOR4_X2__A3_c2 VSS N_A3_M1_g 8.04354e-17
C_x_PM_NOR4_X2__A3_c3 VSS N_A3_M5_g 4.7e-17
R_x_PM_NOR4_X2__A3_r4 x_PM_NOR4_X2__A3_18 x_PM_NOR4_X2__A3_14 4.74714
R_x_PM_NOR4_X2__A3_r5 x_PM_NOR4_X2__A3_17 x_PM_NOR4_X2__A3_14 4.74714
R_x_PM_NOR4_X2__A3_r6 x_PM_NOR4_X2__A3_14 x_PM_NOR4_X2__A3_12 25.0012
R_x_PM_NOR4_X2__A3_r7 x_PM_NOR4_X2__A3_12 A3 0.156071
R_x_PM_NOR4_X2__A3_r8 N_A3_M1_g x_PM_NOR4_X2__A3_18 70.98
R_x_PM_NOR4_X2__A3_r9 N_A3_M5_g x_PM_NOR4_X2__A3_17 42.9
C_x_PM_NOR4_X2__A2_c0 VSS x_PM_NOR4_X2__A2_11 9.40823e-18
C_x_PM_NOR4_X2__A2_c1 VSS x_PM_NOR4_X2__A2_9 7.48156e-17
C_x_PM_NOR4_X2__A2_c2 VSS N_A2_M2_g 7.24567e-17
C_x_PM_NOR4_X2__A2_c3 VSS N_A2_M6_g 5.58007e-17
R_x_PM_NOR4_X2__A2_r4 x_PM_NOR4_X2__A2_18 x_PM_NOR4_X2__A2_11 4.74714
R_x_PM_NOR4_X2__A2_r5 x_PM_NOR4_X2__A2_17 x_PM_NOR4_X2__A2_11 4.74714
R_x_PM_NOR4_X2__A2_r6 x_PM_NOR4_X2__A2_11 x_PM_NOR4_X2__A2_9 25.0012
R_x_PM_NOR4_X2__A2_r7 A2 x_PM_NOR4_X2__A2_9 0.1748
R_x_PM_NOR4_X2__A2_r8 N_A2_M2_g x_PM_NOR4_X2__A2_18 58.5
R_x_PM_NOR4_X2__A2_r9 N_A2_M6_g x_PM_NOR4_X2__A2_17 55.38
C_x_PM_NOR4_X2__A1_c0 VSS x_PM_NOR4_X2__A1_18 1.20639e-17
C_x_PM_NOR4_X2__A1_c1 VSS x_PM_NOR4_X2__A1_9 8.8423e-17
C_x_PM_NOR4_X2__A1_c2 VSS N_A1_M3_g 7.69685e-17
C_x_PM_NOR4_X2__A1_c3 VSS N_A1_M7_g 5.68099e-17
R_x_PM_NOR4_X2__A1_r4 x_PM_NOR4_X2__A1_18 x_PM_NOR4_X2__A1_11 3.38
R_x_PM_NOR4_X2__A1_r5 x_PM_NOR4_X2__A1_11 x_PM_NOR4_X2__A1_9 25.0012
R_x_PM_NOR4_X2__A1_r6 A1 x_PM_NOR4_X2__A1_9 0.198636
R_x_PM_NOR4_X2__A1_r7 x_PM_NOR4_X2__A1_18 x_PM_NOR4_X2__A1_5 1.95
R_x_PM_NOR4_X2__A1_r8 N_A1_M3_g x_PM_NOR4_X2__A1_5 58.5
R_x_PM_NOR4_X2__A1_r9 x_PM_NOR4_X2__A1_18 x_PM_NOR4_X2__A1_VSS 1.95
R_x_PM_NOR4_X2__A1_r10 N_A1_M7_g x_PM_NOR4_X2__A1_VSS 55.38
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
