module singlepath (a0, s31);
input a0;
output s31;
wire w312, w311, w302, w301, c30, w291, s27, c28, c27, s26, w262, s25, c26, w261, w252, w242, w241, s23, c24, w232, w231, w251, c23, c25, w221, c22, w212, w192, s19, w191, s18, w182, c18, w172, w292, w171, w162, w161, w152, w151, w51, s6, s21, s10, w22, w282, w62, c29, s3, c31, c16, c4, w61, c5, s24, w32, w00, s29, w21, s5, w222, w41, s11, w272, w201, c6, c1, w03, s2, w141, w52, w42, w11, w111, s28, w181, w71, s12, s1, s15, w12, w211, c20, c3, s17, c17, w72, c8, s20, s7, w122, c21, w81, s16, w31, w82, w202, c2, c9, s8, w91, s30, w92, c10, c14, s9, c19, s4, w102, w121, c11, w112, w281, w02, c12, w271, w132, c7, c13, s14, w131, s13, w142, s22, w101, c15, Vcc, gnd;
and g0(w00, a0, Vcc);
and g2(w02, a0, Vcc);
or g3(c1, w00, gnd, gnd);
xor g4(w03, a0, gnd);
and ag1(w11, c1, Vcc);
and ag2(w12, c1, Vcc);
or ag3(c2, w12, gnd, gnd);
xor ag5(s1, c1, gnd);
and bg1(w21, c2, Vcc);
and bg2(w22, c2, Vcc);
or bg3(c3, w22, gnd, gnd);
xor bg5(s2, c2, gnd);
and cg1(w31, c3, Vcc);
and cg2(w32, c3, Vcc);
or cg3(c4, w32, gnd, gnd);
xor cg5(s3, c3, gnd);
and dg1(w41, c4, Vcc);
and dg2(w42, c4, Vcc);
or dg3(c5, w42, gnd, gnd);
xor dg5(s4, c4, gnd);
and eg1(w51, c5, Vcc);
and eg2(w52, c5, Vcc);
or eg3(c6, w52, gnd, gnd);
xor eg5(s5, c5, gnd);
and fg1(w61, c6, Vcc);
and fg2(w62, c6, Vcc);
or fg3(c7, w62, gnd, gnd);
xor fg5(s6, c6, gnd);
and gg1(w71, c7, Vcc);
and gg2(w72, c7, Vcc);
or gg3(c8, w72, gnd, gnd);
xor gg5(s7, c7, gnd);
and hg1(w81, c8, Vcc);
and hg2(w82, c8, Vcc);
or hg3(c9, w82, gnd, gnd);
xor hg5(s8, c8, gnd);
and ig1(w91, c9, Vcc);
and ig2(w92, c9, Vcc);
or ig3(c10, w92, gnd, gnd);
xor ig5(s9, c9, gnd);
and jg1(w101, c10, Vcc);
and jg2(w102, c10, Vcc);
or jg3(c11, w102, gnd, gnd);
xor jg5(s10, c10, gnd);
and kg1(w111, c11, Vcc);
and kg2(w112, c11, Vcc);
or kg3(c12, w112, gnd, gnd);
xor kg5(s11, c11, gnd);
and lg1(w121, c12, Vcc);
and lg2(w122, c12, Vcc);
or lg3(c13, w122, gnd, gnd);
xor lg5(s12, c12, gnd);
and mg1(w131, c13, Vcc);
and mg2(w132, c13, Vcc);
or mg3(c14, w132, gnd, gnd);
xor mg5(s13, c13, gnd);
and ng1(w141, c14, Vcc);
and ng2(w142, c14, Vcc);
or ng3(c15, w142, gnd, gnd);
xor ng5(s14, c14, gnd);
and og1(w151, c15, Vcc);
and og2(w152, c15, Vcc);
or og3(c16, w152, gnd, gnd);
xor og5(s15, c15, gnd);
and pg1(w161, c16, Vcc);
and pg2(w162, c16, Vcc);
or pg3(c17, w162, gnd, gnd);
xor pg5(s16, c16, gnd);
and qg1(w171, c17, Vcc);
and qg2(w172, c17, Vcc);
or qg3(c18, w172, gnd, gnd);
xor qg5(s17, c17, gnd);
and rg1(w181, c18, Vcc);
and rg2(w182, c18, Vcc);
or rg3(c19, w182, gnd, gnd);
xor rg5(s18, c18, gnd);
and sg1(w191, c19, Vcc);
and sg2(w192, c19, Vcc);
or sg3(c20, w192, gnd, gnd);
xor sg5(s19, c19, gnd);
and tg1(w201, c20, Vcc);
and tg2(w202, c20, Vcc);
or tg3(c21, w202, gnd, gnd);
xor tg5(s20, c20, gnd);
and ug1(w211, c21, Vcc);
and ug2(w212, c21, Vcc);
or ug3(c22, w212, gnd, gnd);
xor ug5(s21, c21, gnd);
and vg1(w221, c22, Vcc);
and vg2(w222, c22, Vcc);
or vg3(c23, w222, gnd, gnd);
xor vg5(s22, c22, gnd);
and wg1(w231, c23, Vcc);
and wg2(w232, c23, Vcc);
or wg3(c24, w232, gnd, gnd);
xor wg5(s23, c23, gnd);
and yg1(w241, c24, Vcc);
and yg2(w242, c24, Vcc);
or yg3(c25, w242, gnd, gnd);
xor yg5(s24, c24, gnd);
and zg1(w251, c25, Vcc);
and zg2(w252, c25, Vcc);
or zg3(c26, w252, gnd, gnd);
xor zg5(s25, c25, gnd);
and g1a(w261, c26, Vcc);
and g2a(w262, c26, Vcc);
or g3a(c27, w262, gnd, gnd);
xor g5a(s26, c26, gnd);
and g1b(w271, c27, Vcc);
and g2b(w272, c27, Vcc);
or g3b(c28, w272, gnd, gnd);
xor g5b(s27, c27, gnd);
and g1c(w281, c28, Vcc);
and g2c(w282, c28, Vcc);
or g3c(c29, w282, gnd, gnd);
xor g5c(s28, c28, gnd);
and g1d(w291, c29, Vcc);
and g2d(w292, c29, Vcc);
or g3d(c30, w292, gnd, gnd);
xor g5d(s29, c29, gnd);
and g1e(w301, c30, Vcc);
and g2e(w302, c30, Vcc);
or g3e(c31, w302, gnd, gnd);
xor g5e(s30, c30, gnd);
and g1f(w311, c31, Vcc);
and g2f(w312, c31, Vcc);
xor g5f(s31, c31, gnd);

endmodule
