.SUBCKT and2 A1 A2 VDD VSS ZN
M_M3 N_3_M0_d N_A1_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.135000U  AS=0.014175P AD=0.018900P PS=0.480000U PD=0.550000U
M_M4 N_VDD_M1_d N_A2_M1_g N_3_M0_d VDD PMOS_VTL L=0.050U W=0.135000U  AS=0.018900P AD=0.028350P PS=0.550000U PD=0.820000U
M_M5 N_ZN_M2_d N_3_M2_g N_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.270000U  AS=0.028350P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 7 N_A1_M3_g N_3_M3_s VSS NMOS_VTL L=0.050U W=0.130000U  AS=0.013650P AD=0.018200P PS=0.470000U PD=0.540000U
M_M1 N_VSS_M4_d N_A2_M4_g 7 VSS NMOS_VTL L=0.050U W=0.130000U  AS=0.018200P AD=0.021700P PS=0.540000U PD=0.640000U
M_M2 N_ZN_M5_d N_3_M5_g N_VSS_M4_d VSS NMOS_VTL L=0.050U W=0.180000U  AS=0.021700P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_AND2_X2__VSS_c0 VSS x_PM_AND2_X2__VSS_12 3.57664e-17
C_x_PM_AND2_X2__VSS_c1 VSS N_VSS_M4_d 3.3282e-17
C_x_PM_AND2_X2__VSS_c2 VSS x_PM_AND2_X2__VSS_2 5.54251e-17
R_x_PM_AND2_X2__VSS_r3 x_PM_AND2_X2__VSS_12 x_PM_AND2_X2__VSS_6 0.145286
R_x_PM_AND2_X2__VSS_r4 N_VSS_M4_d x_PM_AND2_X2__VSS_6 0.420714
R_x_PM_AND2_X2__VSS_r5 x_PM_AND2_X2__VSS_12 x_PM_AND2_X2__VSS_2 0.0731438
R_x_PM_AND2_X2__VSS_r6 VSS x_PM_AND2_X2__VSS_2 0.0782353
C_x_PM_AND2_X2__VDD_c0 VSS x_PM_AND2_X2__VDD_17 4.42012e-17
C_x_PM_AND2_X2__VDD_c1 VSS N_VDD_M1_d 3.53236e-17
C_x_PM_AND2_X2__VDD_c2 VSS x_PM_AND2_X2__VDD_8 1.07001e-17
C_x_PM_AND2_X2__VDD_c3 VSS x_PM_AND2_X2__VDD_7 3.2606e-17
C_x_PM_AND2_X2__VDD_c4 VSS N_VDD_M0_s 1.42739e-17
R_x_PM_AND2_X2__VDD_r5 x_PM_AND2_X2__VDD_17 x_PM_AND2_X2__VDD_11 0.145286
R_x_PM_AND2_X2__VDD_r6 N_VDD_M1_d x_PM_AND2_X2__VDD_11 0.420714
R_x_PM_AND2_X2__VDD_r7 VDD x_PM_AND2_X2__VDD_8 0.603529
R_x_PM_AND2_X2__VDD_r8 x_PM_AND2_X2__VDD_17 x_PM_AND2_X2__VDD_7 0.0731438
R_x_PM_AND2_X2__VDD_r9 VDD x_PM_AND2_X2__VDD_7 0.0894118
R_x_PM_AND2_X2__VDD_r10 x_PM_AND2_X2__VDD_8 x_PM_AND2_X2__VDD_3 0.264221
R_x_PM_AND2_X2__VDD_r11 N_VDD_M0_s x_PM_AND2_X2__VDD_3 0.420714
C_x_PM_AND2_X2__3_c0 VSS x_PM_AND2_X2__3_33 1.13133e-17
C_x_PM_AND2_X2__3_c1 VSS x_PM_AND2_X2__3_30 1.00152e-17
C_x_PM_AND2_X2__3_c2 VSS x_PM_AND2_X2__3_29 9.34287e-17
C_x_PM_AND2_X2__3_c3 VSS x_PM_AND2_X2__3_26 1.87365e-17
C_x_PM_AND2_X2__3_c4 VSS x_PM_AND2_X2__3_22 8.60574e-18
C_x_PM_AND2_X2__3_c5 VSS x_PM_AND2_X2__3_21 4.03179e-17
C_x_PM_AND2_X2__3_c6 VSS N_3_M0_d 3.31237e-17
C_x_PM_AND2_X2__3_c7 VSS x_PM_AND2_X2__3_16 5.73522e-18
C_x_PM_AND2_X2__3_c8 VSS x_PM_AND2_X2__3_15 6.02033e-17
C_x_PM_AND2_X2__3_c9 VSS N_3_M3_s 2.55776e-17
C_x_PM_AND2_X2__3_c10 VSS N_3_M2_g 9.71074e-17
C_x_PM_AND2_X2__3_c11 VSS N_3_M5_g 3.53623e-17
R_x_PM_AND2_X2__3_r12 x_PM_AND2_X2__3_33 x_PM_AND2_X2__3_31 3.38
R_x_PM_AND2_X2__3_r13 x_PM_AND2_X2__3_29 x_PM_AND2_X2__3_30 2.93143
R_x_PM_AND2_X2__3_r14 x_PM_AND2_X2__3_31 x_PM_AND2_X2__3_26 25.0012
R_x_PM_AND2_X2__3_r15 x_PM_AND2_X2__3_30 x_PM_AND2_X2__3_24 0.232321
R_x_PM_AND2_X2__3_r16 x_PM_AND2_X2__3_26 x_PM_AND2_X2__3_24 0.0542857
R_x_PM_AND2_X2__3_r17 x_PM_AND2_X2__3_26 x_PM_AND2_X2__3_23 0.22619
R_x_PM_AND2_X2__3_r18 x_PM_AND2_X2__3_29 x_PM_AND2_X2__3_21 0.212317
R_x_PM_AND2_X2__3_r19 x_PM_AND2_X2__3_22 x_PM_AND2_X2__3_21 0.76
R_x_PM_AND2_X2__3_r20 x_PM_AND2_X2__3_22 x_PM_AND2_X2__3_17 0.212317
R_x_PM_AND2_X2__3_r21 N_3_M0_d x_PM_AND2_X2__3_17 0.393571
R_x_PM_AND2_X2__3_r22 x_PM_AND2_X2__3_23 x_PM_AND2_X2__3_15 0.223553
R_x_PM_AND2_X2__3_r23 x_PM_AND2_X2__3_16 x_PM_AND2_X2__3_15 1.79143
R_x_PM_AND2_X2__3_r24 x_PM_AND2_X2__3_16 x_PM_AND2_X2__3_11 0.212317
R_x_PM_AND2_X2__3_r25 N_3_M3_s x_PM_AND2_X2__3_11 0.420714
R_x_PM_AND2_X2__3_r26 x_PM_AND2_X2__3_33 x_PM_AND2_X2__3_5 1.95
R_x_PM_AND2_X2__3_r27 N_3_M2_g x_PM_AND2_X2__3_5 105.3
R_x_PM_AND2_X2__3_r28 x_PM_AND2_X2__3_33 x_PM_AND2_X2__3_VSS 1.95
R_x_PM_AND2_X2__3_r29 N_3_M5_g x_PM_AND2_X2__3_VSS 27.3
C_x_PM_AND2_X2__A1_c0 VSS x_PM_AND2_X2__A1_13 7.02743e-18
C_x_PM_AND2_X2__A1_c1 VSS A1 1.56682e-17
C_x_PM_AND2_X2__A1_c2 VSS N_A1_M0_g 6.18939e-17
C_x_PM_AND2_X2__A1_c3 VSS N_A1_M3_g 5.49708e-17
R_x_PM_AND2_X2__A1_r4 x_PM_AND2_X2__A1_16 x_PM_AND2_X2__A1_13 4.74714
R_x_PM_AND2_X2__A1_r5 x_PM_AND2_X2__A1_15 x_PM_AND2_X2__A1_13 4.74714
R_x_PM_AND2_X2__A1_r6 x_PM_AND2_X2__A1_13 x_PM_AND2_X2__A1_11 25.0012
R_x_PM_AND2_X2__A1_r7 x_PM_AND2_X2__A1_11 A1 0.158563
R_x_PM_AND2_X2__A1_r8 N_A1_M0_g x_PM_AND2_X2__A1_16 83.85
R_x_PM_AND2_X2__A1_r9 N_A1_M3_g x_PM_AND2_X2__A1_15 63.18
C_x_PM_AND2_X2__A2_c0 VSS x_PM_AND2_X2__A2_14 8.64377e-18
C_x_PM_AND2_X2__A2_c1 VSS x_PM_AND2_X2__A2_12 4.37781e-17
C_x_PM_AND2_X2__A2_c2 VSS N_A2_M1_g 5.57959e-17
C_x_PM_AND2_X2__A2_c3 VSS N_A2_M4_g 7.00537e-17
R_x_PM_AND2_X2__A2_r4 x_PM_AND2_X2__A2_18 x_PM_AND2_X2__A2_14 4.7687
R_x_PM_AND2_X2__A2_r5 x_PM_AND2_X2__A2_17 x_PM_AND2_X2__A2_14 4.7687
R_x_PM_AND2_X2__A2_r6 x_PM_AND2_X2__A2_14 x_PM_AND2_X2__A2_12 25.0012
R_x_PM_AND2_X2__A2_r7 x_PM_AND2_X2__A2_12 A2 0.169643
R_x_PM_AND2_X2__A2_r8 N_A2_M1_g x_PM_AND2_X2__A2_18 62.01
R_x_PM_AND2_X2__A2_r9 N_A2_M4_g x_PM_AND2_X2__A2_17 85.02
C_x_PM_AND2_X2__ZN_c0 VSS N_ZN_M5_d 2.60988e-17
C_x_PM_AND2_X2__ZN_c1 VSS ZN 7.63258e-17
C_x_PM_AND2_X2__ZN_c2 VSS N_ZN_M2_d 5.16564e-17
C_x_PM_AND2_X2__ZN_c3 VSS x_PM_AND2_X2__ZN_3 6.61381e-18
R_x_PM_AND2_X2__ZN_r4 ZN x_PM_AND2_X2__ZN_8 1.87286
R_x_PM_AND2_X2__ZN_r5 x_PM_AND2_X2__ZN_7 N_ZN_M5_d 0.30478
R_x_PM_AND2_X2__ZN_r6 ZN x_PM_AND2_X2__ZN_7 1.60143
R_x_PM_AND2_X2__ZN_r7 x_PM_AND2_X2__ZN_8 x_PM_AND2_X2__ZN_3 0.20978
R_x_PM_AND2_X2__ZN_r8 N_ZN_M2_d x_PM_AND2_X2__ZN_3 0.686111
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
