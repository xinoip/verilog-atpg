
module c3540_tb();



reg N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
      N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
      N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
      N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
      N303,N311,N317,N322,N326,N329,N330,N343,N349,N350;

wire N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
       N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
       N5360,N5361;
	
	 
c3540 c0(N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
		  N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
		  N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
		  N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
		  N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,
		  N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
		  N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
		  N5360,N5361);	
	 
reg [49:0] test_vectors[0:9];	
reg [21:0] out_vectors[0:9];	

integer k;
			 
initial
	begin

	$readmemb("c3540_input_data.txt", test_vectors);
	
	end
	
initial
	begin
	
	for(k = 0; k < 10; k = k + 1)
		begin		
		#10
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
      N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
      N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
      N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
      N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = test_vectors[k];
			
		#1
		out_vectors[k] = {N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
       N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
       N5360,N5361};
		 
		$display("output%d: %h\n", k, out_vectors[k]);
		
		end
		
		$writememb("c3540_in_data.txt", test_vectors);
		$writememb("c3540_out_data.txt", out_vectors);
	
	end



endmodule
