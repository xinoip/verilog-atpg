.SUBCKT nor8 A1 A2 A3 A4 A5 A6 A7 A8 VDD VSS ZN
************************************************NOR4_X2********************************************
M_M4 8 N_A4_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.650000U AS=0.068250P AD=0.091000P PS=1.510000U PD=1.580000U
M_M5 9 N_A3_M1_g 8 VDD PMOS_VTL L=0.050U W=0.650000U AS=0.091000P AD=0.091000P PS=1.580000U PD=1.580000U
M_M6 10 N_A2_M2_g 9 VDD PMOS_VTL L=0.050U W=0.650000U AS=0.091000P AD=0.091000P PS=1.580000U PD=1.580000U
M_M7 N_Zalp1_M3_d N_A1_M3_g 10 VDD PMOS_VTL L=0.050U W=0.650000U AS=0.091000P AD=0.068250P PS=1.580000U PD=1.510000U
M_M0 N_Zalp1_M4_d N_A4_M4_g N_VSS_M4_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M_M1 N_VSS_M5_d N_A3_M5_g N_Zalp1_M4_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M_M2 N_Zalp1_M6_d N_A2_M6_g N_VSS_M5_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M_M3 N_VSS_M7_d N_A1_M7_g N_Zalp1_M6_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_NOR4_X2__VSS_c0 VSS VSS 2.64443e-18
C_x_PM_NOR4_X2__VSS_c1 VSS N_VSS_M7_d 1.30717e-17
C_x_PM_NOR4_X2__VSS_c2 VSS x_PM_NOR4_X2__VSS_14 5.3438e-17
C_x_PM_NOR4_X2__VSS_c3 VSS N_VSS_M5_d 2.04204e-17
C_x_PM_NOR4_X2__VSS_c4 VSS x_PM_NOR4_X2__VSS_9 1.06295e-17
C_x_PM_NOR4_X2__VSS_c5 VSS x_PM_NOR4_X2__VSS_8 3.88904e-17
C_x_PM_NOR4_X2__VSS_c6 VSS N_VSS_M4_s 1.0831e-17
R_x_PM_NOR4_X2__VSS_r7 N_VSS_M7_d x_PM_NOR4_X2__VSS_16 0.230714
R_x_PM_NOR4_X2__VSS_r8 VSS x_PM_NOR4_X2__VSS_15 0.0731438
R_x_PM_NOR4_X2__VSS_r9 x_PM_NOR4_X2__VSS_16 x_PM_NOR4_X2__VSS_14 0.264221
R_x_PM_NOR4_X2__VSS_r10 x_PM_NOR4_X2__VSS_15 x_PM_NOR4_X2__VSS_14 0.681765
R_x_PM_NOR4_X2__VSS_r11 VSS x_PM_NOR4_X2__VSS_10 0.145286
R_x_PM_NOR4_X2__VSS_r12 N_VSS_M5_d x_PM_NOR4_X2__VSS_10 0.230714
R_x_PM_NOR4_X2__VSS_r13 VSS x_PM_NOR4_X2__VSS_8 0.0731438
R_x_PM_NOR4_X2__VSS_r14 x_PM_NOR4_X2__VSS_9 x_PM_NOR4_X2__VSS_8 0.692941
R_x_PM_NOR4_X2__VSS_r15 x_PM_NOR4_X2__VSS_9 x_PM_NOR4_X2__VSS_4 0.264221
R_x_PM_NOR4_X2__VSS_r16 N_VSS_M4_s x_PM_NOR4_X2__VSS_4 0.230714
C_x_PM_NOR4_X2__VDD_c0 VSS VDD 7.40695e-17
C_x_PM_NOR4_X2__VDD_c1 VSS N_VDD_M0_s 2.4691e-17
C_x_PM_NOR4_X2__VDD_c2 VSS x_PM_NOR4_X2__VDD_2 1.06862e-17
R_x_PM_NOR4_X2__VDD_r3 VDD x_PM_NOR4_X2__VDD_2 0.0689273
R_x_PM_NOR4_X2__VDD_r4 N_VDD_M0_s x_PM_NOR4_X2__VDD_2 0.230714
C_x_PM_NOR4_X2__A4_c0 VSS x_PM_NOR4_X2__A4_14 7.18659e-18
C_x_PM_NOR4_X2__A4_c1 VSS x_PM_NOR4_X2__A4_12 3.56769e-17
C_x_PM_NOR4_X2__A4_c2 VSS N_A4_M0_g 7.98018e-17
C_x_PM_NOR4_X2__A4_c3 VSS N_A4_M4_g 4.23053e-17
R_x_PM_NOR4_X2__A4_r4 x_PM_NOR4_X2__A4_18 x_PM_NOR4_X2__A4_14 4.74714
R_x_PM_NOR4_X2__A4_r5 x_PM_NOR4_X2__A4_17 x_PM_NOR4_X2__A4_14 4.74714
R_x_PM_NOR4_X2__A4_r6 x_PM_NOR4_X2__A4_14 x_PM_NOR4_X2__A4_12 25.0012
R_x_PM_NOR4_X2__A4_r7 x_PM_NOR4_X2__A4_12 A4 0.156071
R_x_PM_NOR4_X2__A4_r8 N_A4_M0_g x_PM_NOR4_X2__A4_18 70.98
R_x_PM_NOR4_X2__A4_r9 N_A4_M4_g x_PM_NOR4_X2__A4_17 42.9
C_x_PM_NOR4_X2__Zalp1_c0 VSS x_PM_NOR4_X2__Zalp1_27 1.32309e-17
C_x_PM_NOR4_X2__Zalp1_c1 VSS x_PM_NOR4_X2__Zalp1_26 2.32902e-17
C_x_PM_NOR4_X2__Zalp1_c2 VSS x_PM_NOR4_X2__Zalp1_23 4.60612e-17
C_x_PM_NOR4_X2__Zalp1_c3 VSS N_Zalp1_M3_d 2.50235e-17
C_x_PM_NOR4_X2__Zalp1_c4 VSS x_PM_NOR4_X2__Zalp1_18 3.46798e-18
C_x_PM_NOR4_X2__Zalp1_c5 VSS x_PM_NOR4_X2__Zalp1_16 2.65091e-17
C_x_PM_NOR4_X2__Zalp1_c6 VSS N_Zalp1_M6_d 2.42211e-17
C_x_PM_NOR4_X2__Zalp1_c7 VSS x_PM_NOR4_X2__Zalp1_11 2.27649e-17
C_x_PM_NOR4_X2__Zalp1_c8 VSS x_PM_NOR4_X2__Zalp1_10 1.9661e-17
C_x_PM_NOR4_X2__Zalp1_c9 VSS x_PM_NOR4_X2__Zalp1_9 1.62159e-17
C_x_PM_NOR4_X2__Zalp1_c10 VSS N_Zalp1_M4_d 2.33665e-17
R_x_PM_NOR4_X2__Zalp1_r11 x_PM_NOR4_X2__Zalp1_26 Zalp1 0.189936
R_x_PM_NOR4_X2__Zalp1_r12 x_PM_NOR4_X2__Zalp1_23 x_PM_NOR4_X2__Zalp1_22 1.65571
R_x_PM_NOR4_X2__Zalp1_r13 x_PM_NOR4_X2__Zalp1_23 x_PM_NOR4_X2__Zalp1_18 0.192227
R_x_PM_NOR4_X2__Zalp1_r14 N_Zalp1_M3_d x_PM_NOR4_X2__Zalp1_18 0.861333
R_x_PM_NOR4_X2__Zalp1_r15 x_PM_NOR4_X2__Zalp1_27 x_PM_NOR4_X2__Zalp1_17 0.113465
R_x_PM_NOR4_X2__Zalp1_r16 x_PM_NOR4_X2__Zalp1_22 x_PM_NOR4_X2__Zalp1_16 0.212317
R_x_PM_NOR4_X2__Zalp1_r17 x_PM_NOR4_X2__Zalp1_17 x_PM_NOR4_X2__Zalp1_16 0.705714
R_x_PM_NOR4_X2__Zalp1_r18 x_PM_NOR4_X2__Zalp1_27 x_PM_NOR4_X2__Zalp1_12 0.0883294
R_x_PM_NOR4_X2__Zalp1_r19 N_Zalp1_M6_d x_PM_NOR4_X2__Zalp1_12 0.257857
R_x_PM_NOR4_X2__Zalp1_r20 Zalp1 x_PM_NOR4_X2__Zalp1_11 0.095
R_x_PM_NOR4_X2__Zalp1_r21 x_PM_NOR4_X2__Zalp1_27 x_PM_NOR4_X2__Zalp1_10 0.113465
R_x_PM_NOR4_X2__Zalp1_r22 x_PM_NOR4_X2__Zalp1_11 x_PM_NOR4_X2__Zalp1_10 0.257857
R_x_PM_NOR4_X2__Zalp1_r23 x_PM_NOR4_X2__Zalp1_9 x_PM_NOR4_X2__Zalp1_26 0.732857
R_x_PM_NOR4_X2__Zalp1_r24 x_PM_NOR4_X2__Zalp1_9 x_PM_NOR4_X2__Zalp1_4 0.212317
R_x_PM_NOR4_X2__Zalp1_r25 N_Zalp1_M4_d x_PM_NOR4_X2__Zalp1_4 0.257857
C_x_PM_NOR4_X2__A3_c0 VSS x_PM_NOR4_X2__A3_14 8.988e-18
C_x_PM_NOR4_X2__A3_c1 VSS x_PM_NOR4_X2__A3_12 6.21612e-17
C_x_PM_NOR4_X2__A3_c2 VSS N_A3_M1_g 8.04354e-17
C_x_PM_NOR4_X2__A3_c3 VSS N_A3_M5_g 4.7e-17
R_x_PM_NOR4_X2__A3_r4 x_PM_NOR4_X2__A3_18 x_PM_NOR4_X2__A3_14 4.74714
R_x_PM_NOR4_X2__A3_r5 x_PM_NOR4_X2__A3_17 x_PM_NOR4_X2__A3_14 4.74714
R_x_PM_NOR4_X2__A3_r6 x_PM_NOR4_X2__A3_14 x_PM_NOR4_X2__A3_12 25.0012
R_x_PM_NOR4_X2__A3_r7 x_PM_NOR4_X2__A3_12 A3 0.156071
R_x_PM_NOR4_X2__A3_r8 N_A3_M1_g x_PM_NOR4_X2__A3_18 70.98
R_x_PM_NOR4_X2__A3_r9 N_A3_M5_g x_PM_NOR4_X2__A3_17 42.9
C_x_PM_NOR4_X2__A2_c0 VSS x_PM_NOR4_X2__A2_11 9.40823e-18
C_x_PM_NOR4_X2__A2_c1 VSS x_PM_NOR4_X2__A2_9 7.48156e-17
C_x_PM_NOR4_X2__A2_c2 VSS N_A2_M2_g 7.24567e-17
C_x_PM_NOR4_X2__A2_c3 VSS N_A2_M6_g 5.58007e-17
R_x_PM_NOR4_X2__A2_r4 x_PM_NOR4_X2__A2_18 x_PM_NOR4_X2__A2_11 4.74714
R_x_PM_NOR4_X2__A2_r5 x_PM_NOR4_X2__A2_17 x_PM_NOR4_X2__A2_11 4.74714
R_x_PM_NOR4_X2__A2_r6 x_PM_NOR4_X2__A2_11 x_PM_NOR4_X2__A2_9 25.0012
R_x_PM_NOR4_X2__A2_r7 A2 x_PM_NOR4_X2__A2_9 0.1748
R_x_PM_NOR4_X2__A2_r8 N_A2_M2_g x_PM_NOR4_X2__A2_18 58.5
R_x_PM_NOR4_X2__A2_r9 N_A2_M6_g x_PM_NOR4_X2__A2_17 55.38
C_x_PM_NOR4_X2__A1_c0 VSS x_PM_NOR4_X2__A1_18 1.20639e-17
C_x_PM_NOR4_X2__A1_c1 VSS x_PM_NOR4_X2__A1_9 8.8423e-17
C_x_PM_NOR4_X2__A1_c2 VSS N_A1_M3_g 7.69685e-17
C_x_PM_NOR4_X2__A1_c3 VSS N_A1_M7_g 5.68099e-17
R_x_PM_NOR4_X2__A1_r4 x_PM_NOR4_X2__A1_18 x_PM_NOR4_X2__A1_11 3.38
R_x_PM_NOR4_X2__A1_r5 x_PM_NOR4_X2__A1_11 x_PM_NOR4_X2__A1_9 25.0012
R_x_PM_NOR4_X2__A1_r6 A1 x_PM_NOR4_X2__A1_9 0.198636
R_x_PM_NOR4_X2__A1_r7 x_PM_NOR4_X2__A1_18 x_PM_NOR4_X2__A1_5 1.95
R_x_PM_NOR4_X2__A1_r8 N_A1_M3_g x_PM_NOR4_X2__A1_5 58.5
R_x_PM_NOR4_X2__A1_r9 x_PM_NOR4_X2__A1_18 x_PM_NOR4_X2__A1_VSS 1.95
R_x_PM_NOR4_X2__A1_r10 N_A1_M7_g x_PM_NOR4_X2__A1_VSS 55.38
***************************************************NOR4_X2***********************************************************
M2_M4 82 N2_A8_M0_g N2_VDD_M0_s VDD PMOS_VTL W=0.650000U AS=0.068250P AD=0.091000P PS=1.510000U PD=1.580000U
M2_M5 92 N2_A7_M1_g 82 VDD PMOS_VTL W=0.650000U AS=0.091000P AD=0.091000P PS=1.580000U PD=1.580000U
M2_M6 102 N2_A6_M2_g 92 VDD PMOS_VTL W=0.650000U AS=0.091000P AD=0.091000P PS=1.580000U PD=1.580000U
M2_M7 N2_Zalp2_M3_d N2_A5_M3_g 102 VDD PMOS_VTL W=0.650000U AS=0.091000P AD=0.068250P PS=1.580000U PD=1.510000U
M2_M0 N2_Zalp2_M4_d N2_A8_M4_g N2_VSS_M4_s VSS NMOS_VTL W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M2_M1 N2_VSS_M5_d N2_A7_M5_g N2_Zalp2_M4_d VSS NMOS_VTL W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M2_M2 N2_Zalp2_M6_d N2_A6_M6_g N2_VSS_M5_d VSS NMOS_VTL W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M2_M3 N2_VSS_M7_d N2_A5_M7_g N2_Zalp2_M6_d VSS NMOS_VTL W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x2_PM2_NOR4_X2__VSS_c0 VSS VSS 2.64443e-18
C_x2_PM2_NOR4_X2__VSS_c1 VSS N2_VSS_M7_d 1.30717e-17
C_x2_PM2_NOR4_X2__VSS_c2 VSS x2_PM2_NOR4_X2__VSS_14 5.3438e-17
C_x2_PM2_NOR4_X2__VSS_c3 VSS N2_VSS_M5_d 2.04204e-17
C_x2_PM2_NOR4_X2__VSS_c4 VSS x2_PM2_NOR4_X2__VSS_9 1.06295e-17
C_x2_PM2_NOR4_X2__VSS_c5 VSS x2_PM2_NOR4_X2__VSS_8 3.88904e-17
C_x2_PM2_NOR4_X2__VSS_c6 VSS N2_VSS_M4_s 1.0831e-17
R_x2_PM2_NOR4_X2__VSS_r7 N2_VSS_M7_d x2_PM2_NOR4_X2__VSS_16 0.230714
R_x2_PM2_NOR4_X2__VSS_r8 VSS x2_PM2_NOR4_X2__VSS_15 0.0731438
R_x2_PM2_NOR4_X2__VSS_r9 x2_PM2_NOR4_X2__VSS_16 x2_PM2_NOR4_X2__VSS_14 0.264221
R_x2_PM2_NOR4_X2__VSS_r10 x2_PM2_NOR4_X2__VSS_15 x2_PM2_NOR4_X2__VSS_14 0.681765
R_x2_PM2_NOR4_X2__VSS_r11 VSS x2_PM2_NOR4_X2__VSS_10 0.145286
R_x2_PM2_NOR4_X2__VSS_r12 N2_VSS_M5_d x2_PM2_NOR4_X2__VSS_10 0.230714
R_x2_PM2_NOR4_X2__VSS_r13 VSS x2_PM2_NOR4_X2__VSS_8 0.0731438
R_x2_PM2_NOR4_X2__VSS_r14 x2_PM2_NOR4_X2__VSS_9 x2_PM2_NOR4_X2__VSS_8 0.692941
R_x2_PM2_NOR4_X2__VSS_r15 x2_PM2_NOR4_X2__VSS_9 x2_PM2_NOR4_X2__VSS_4 0.264221
R_x2_PM2_NOR4_X2__VSS_r16 N2_VSS_M4_s x2_PM2_NOR4_X2__VSS_4 0.230714
C_x2_PM2_NOR4_X2__VDD_c0 VSS VDD 7.40695e-17
C_x2_PM2_NOR4_X2__VDD_c1 VSS N2_VDD_M0_s 2.4691e-17
C_x2_PM2_NOR4_X2__VDD_c2 VSS x2_PM2_NOR4_X2__VDD_2 1.06862e-17
R_x2_PM2_NOR4_X2__VDD_r3 VDD x2_PM2_NOR4_X2__VDD_2 0.0689273
R_x2_PM2_NOR4_X2__VDD_r4 N2_VDD_M0_s x2_PM2_NOR4_X2__VDD_2 0.230714
C_x2_PM2_NOR4_X2__A8_c0 VSS x2_PM2_NOR4_X2__A8_14 7.18659e-18
C_x2_PM2_NOR4_X2__A8_c1 VSS x2_PM2_NOR4_X2__A8_12 3.56769e-17
C_x2_PM2_NOR4_X2__A8_c2 VSS N2_A8_M0_g 7.98018e-17
C_x2_PM2_NOR4_X2__A8_c3 VSS N2_A8_M4_g 4.23053e-17
R_x2_PM2_NOR4_X2__A8_r4 x2_PM2_NOR4_X2__A8_18 x2_PM2_NOR4_X2__A8_14 4.74714
R_x2_PM2_NOR4_X2__A8_r5 x2_PM2_NOR4_X2__A8_17 x2_PM2_NOR4_X2__A8_14 4.74714
R_x2_PM2_NOR4_X2__A8_r6 x2_PM2_NOR4_X2__A8_14 x2_PM2_NOR4_X2__A8_12 25.0012
R_x2_PM2_NOR4_X2__A8_r7 x2_PM2_NOR4_X2__A8_12 A8 0.156071
R_x2_PM2_NOR4_X2__A8_r8 N2_A8_M0_g x2_PM2_NOR4_X2__A8_18 70.98
R_x2_PM2_NOR4_X2__A8_r9 N2_A8_M4_g x2_PM2_NOR4_X2__A8_17 42.9
C_x2_PM2_NOR4_X2__Zalp2_c0 VSS x2_PM2_NOR4_X2__Zalp2_27 1.32309e-17
C_x2_PM2_NOR4_X2__Zalp2_c1 VSS x2_PM2_NOR4_X2__Zalp2_26 2.32902e-17
C_x2_PM2_NOR4_X2__Zalp2_c2 VSS x2_PM2_NOR4_X2__Zalp2_23 4.60612e-17
C_x2_PM2_NOR4_X2__Zalp2_c3 VSS N2_Zalp2_M3_d 2.50235e-17
C_x2_PM2_NOR4_X2__Zalp2_c4 VSS x2_PM2_NOR4_X2__Zalp2_18 3.46798e-18
C_x2_PM2_NOR4_X2__Zalp2_c5 VSS x2_PM2_NOR4_X2__Zalp2_16 2.65091e-17
C_x2_PM2_NOR4_X2__Zalp2_c6 VSS N2_Zalp2_M6_d 2.42211e-17
C_x2_PM2_NOR4_X2__Zalp2_c7 VSS x2_PM2_NOR4_X2__Zalp2_11 2.27649e-17
C_x2_PM2_NOR4_X2__Zalp2_c8 VSS x2_PM2_NOR4_X2__Zalp2_10 1.9661e-17
C_x2_PM2_NOR4_X2__Zalp2_c9 VSS x2_PM2_NOR4_X2__Zalp2_9 1.62159e-17
C_x2_PM2_NOR4_X2__Zalp2_c10 VSS N2_Zalp2_M4_d 2.33665e-17
R_x2_PM2_NOR4_X2__Zalp2_r11 x2_PM2_NOR4_X2__Zalp2_26 Zalp2 0.189936
R_x2_PM2_NOR4_X2__Zalp2_r12 x2_PM2_NOR4_X2__Zalp2_23 x2_PM2_NOR4_X2__Zalp2_22 1.65571
R_x2_PM2_NOR4_X2__Zalp2_r13 x2_PM2_NOR4_X2__Zalp2_23 x2_PM2_NOR4_X2__Zalp2_18 0.192227
R_x2_PM2_NOR4_X2__Zalp2_r14 N2_Zalp2_M3_d x2_PM2_NOR4_X2__Zalp2_18 0.861333
R_x2_PM2_NOR4_X2__Zalp2_r15 x2_PM2_NOR4_X2__Zalp2_27 x2_PM2_NOR4_X2__Zalp2_17 0.113465
R_x2_PM2_NOR4_X2__Zalp2_r16 x2_PM2_NOR4_X2__Zalp2_22 x2_PM2_NOR4_X2__Zalp2_16 0.212317
R_x2_PM2_NOR4_X2__Zalp2_r17 x2_PM2_NOR4_X2__Zalp2_17 x2_PM2_NOR4_X2__Zalp2_16 0.705714
R_x2_PM2_NOR4_X2__Zalp2_r18 x2_PM2_NOR4_X2__Zalp2_27 x2_PM2_NOR4_X2__Zalp2_12 0.0883294
R_x2_PM2_NOR4_X2__Zalp2_r19 N2_Zalp2_M6_d x2_PM2_NOR4_X2__Zalp2_12 0.257857
R_x2_PM2_NOR4_X2__Zalp2_r20 Zalp2 x2_PM2_NOR4_X2__Zalp2_11 0.095
R_x2_PM2_NOR4_X2__Zalp2_r21 x2_PM2_NOR4_X2__Zalp2_27 x2_PM2_NOR4_X2__Zalp2_10 0.113465
R_x2_PM2_NOR4_X2__Zalp2_r22 x2_PM2_NOR4_X2__Zalp2_11 x2_PM2_NOR4_X2__Zalp2_10 0.257857
R_x2_PM2_NOR4_X2__Zalp2_r23 x2_PM2_NOR4_X2__Zalp2_9 x2_PM2_NOR4_X2__Zalp2_26 0.732857
R_x2_PM2_NOR4_X2__Zalp2_r24 x2_PM2_NOR4_X2__Zalp2_9 x2_PM2_NOR4_X2__Zalp2_4 0.212317
R_x2_PM2_NOR4_X2__Zalp2_r25 N2_Zalp2_M4_d x2_PM2_NOR4_X2__Zalp2_4 0.257857
C_x2_PM2_NOR4_X2__A7_c0 VSS x2_PM2_NOR4_X2__A7_14 8.988e-18
C_x2_PM2_NOR4_X2__A7_c1 VSS x2_PM2_NOR4_X2__A7_12 6.21612e-17
C_x2_PM2_NOR4_X2__A7_c2 VSS N2_A7_M1_g 8.04354e-17
C_x2_PM2_NOR4_X2__A7_c3 VSS N2_A7_M5_g 4.7e-17
R_x2_PM2_NOR4_X2__A7_r4 x2_PM2_NOR4_X2__A7_18 x2_PM2_NOR4_X2__A7_14 4.74714
R_x2_PM2_NOR4_X2__A7_r5 x2_PM2_NOR4_X2__A7_17 x2_PM2_NOR4_X2__A7_14 4.74714
R_x2_PM2_NOR4_X2__A7_r6 x2_PM2_NOR4_X2__A7_14 x2_PM2_NOR4_X2__A7_12 25.0012
R_x2_PM2_NOR4_X2__A7_r7 x2_PM2_NOR4_X2__A7_12 A7 0.156071
R_x2_PM2_NOR4_X2__A7_r8 N2_A7_M1_g x2_PM2_NOR4_X2__A7_18 70.98
R_x2_PM2_NOR4_X2__A7_r9 N2_A7_M5_g x2_PM2_NOR4_X2__A7_17 42.9
C_x2_PM2_NOR4_X2__A6_c0 VSS x2_PM2_NOR4_X2__A6_11 9.40823e-18
C_x2_PM2_NOR4_X2__A6_c1 VSS x2_PM2_NOR4_X2__A6_9 7.48156e-17
C_x2_PM2_NOR4_X2__A6_c2 VSS N2_A6_M2_g 7.24567e-17
C_x2_PM2_NOR4_X2__A6_c3 VSS N2_A6_M6_g 5.58007e-17
R_x2_PM2_NOR4_X2__A6_r4 x2_PM2_NOR4_X2__A6_18 x2_PM2_NOR4_X2__A6_11 4.74714
R_x2_PM2_NOR4_X2__A6_r5 x2_PM2_NOR4_X2__A6_17 x2_PM2_NOR4_X2__A6_11 4.74714
R_x2_PM2_NOR4_X2__A6_r6 x2_PM2_NOR4_X2__A6_11 x2_PM2_NOR4_X2__A6_9 25.0012
R_x2_PM2_NOR4_X2__A6_r7 A6 x2_PM2_NOR4_X2__A6_9 0.1748
R_x2_PM2_NOR4_X2__A6_r8 N2_A6_M2_g x2_PM2_NOR4_X2__A6_18 58.5
R_x2_PM2_NOR4_X2__A6_r9 N2_A6_M6_g x2_PM2_NOR4_X2__A6_17 55.38
C_x2_PM2_NOR4_X2__A5_c0 VSS x2_PM2_NOR4_X2__A5_18 1.20639e-17
C_x2_PM2_NOR4_X2__A5_c1 VSS x2_PM2_NOR4_X2__A5_9 8.8423e-17
C_x2_PM2_NOR4_X2__A5_c2 VSS N2_A5_M3_g 7.69685e-17
C_x2_PM2_NOR4_X2__A5_c3 VSS N2_A5_M7_g 5.68099e-17
R_x2_PM2_NOR4_X2__A5_r4 x2_PM2_NOR4_X2__A5_18 x2_PM2_NOR4_X2__A5_11 3.38
R_x2_PM2_NOR4_X2__A5_r5 x2_PM2_NOR4_X2__A5_11 x2_PM2_NOR4_X2__A5_9 25.0012
R_x2_PM2_NOR4_X2__A5_r6 A5 x2_PM2_NOR4_X2__A5_9 0.198636
R_x2_PM2_NOR4_X2__A5_r7 x2_PM2_NOR4_X2__A5_18 x2_PM2_NOR4_X2__A5_5 1.95
R_x2_PM2_NOR4_X2__A5_r8 N2_A5_M3_g x2_PM2_NOR4_X2__A5_5 58.5
R_x2_PM2_NOR4_X2__A5_r9 x2_PM2_NOR4_X2__A5_18 x2_PM2_NOR4_X2__A5_VSS 1.95
R_x2_PM2_NOR4_X2__A5_r10 N2_A5_M7_g x2_PM2_NOR4_X2__A5_VSS 55.38
******************************************************AND2_X2******************************************************
M3_M3 N3_3_M0_d N3_Zalp1_M0_g N3_VDD_M0_s VDD PMOS_VTL W=0.135000U  AS=0.014175P AD=0.018900P PS=0.480000U PD=0.550000U
M3_M4 N3_VDD_M1_d N3_Zalp2_M1_g N3_3_M0_d VDD PMOS_VTL W=0.135000U  AS=0.018900P AD=0.028350P PS=0.550000U PD=0.820000U
M3_M5 N3_ZN3_M2_d N3_3_M2_g N3_VDD_M1_d VDD PMOS_VTL W=0.270000U  AS=0.028350P AD=0.028350P PS=0.820000U PD=0.750000U
M3_M0 73 N3_Zalp1_M3_g N3_3_M3_s VSS NMOS_VTL W=0.130000U  AS=0.013650P AD=0.018200P PS=0.470000U PD=0.540000U
M3_M1 N3_VSS_M4_d N3_Zalp2_M4_g 73 VSS NMOS_VTL W=0.130000U  AS=0.018200P AD=0.021700P PS=0.540000U PD=0.640000U
M3_M2 N3_ZN3_M5_d N3_3_M5_g N3_VSS_M4_d VSS NMOS_VTL W=0.180000U  AS=0.021700P AD=0.018900P PS=0.640000U PD=0.570000U
C_x3_PM_AND2_X2__VSS_c0 VSS x3_PM_AND2_X2__VSS_12 3.57664e-17
C_x3_PM_AND2_X2__VSS_c1 VSS N3_VSS_M4_d 3.3282e-17
C_x3_PM_AND2_X2__VSS_c2 VSS x3_PM_AND2_X2__VSS_2 5.54251e-17
R_x3_PM_AND2_X2__VSS_r3 x3_PM_AND2_X2__VSS_12 x3_PM_AND2_X2__VSS_6 0.145286
R_x3_PM_AND2_X2__VSS_r4 N3_VSS_M4_d x3_PM_AND2_X2__VSS_6 0.420714
R_x3_PM_AND2_X2__VSS_r5 x3_PM_AND2_X2__VSS_12 x3_PM_AND2_X2__VSS_2 0.0731438
R_x3_PM_AND2_X2__VSS_r6 VSS x3_PM_AND2_X2__VSS_2 0.0782353
C_x3_PM_AND2_X2__VDD_c0 VSS x3_PM_AND2_X2__VDD_17 4.42012e-17
C_x3_PM_AND2_X2__VDD_c1 VSS N3_VDD_M1_d 3.53236e-17
C_x3_PM_AND2_X2__VDD_c2 VSS x3_PM_AND2_X2__VDD_8 1.07001e-17
C_x3_PM_AND2_X2__VDD_c3 VSS x3_PM_AND2_X2__VDD_7 3.2606e-17
C_x3_PM_AND2_X2__VDD_c4 VSS N3_VDD_M0_s 1.42739e-17
R_x3_PM_AND2_X2__VDD_r5 x3_PM_AND2_X2__VDD_17 x3_PM_AND2_X2__VDD_11 0.145286
R_x3_PM_AND2_X2__VDD_r6 N3_VDD_M1_d x3_PM_AND2_X2__VDD_11 0.420714
R_x3_PM_AND2_X2__VDD_r7 VDD x3_PM_AND2_X2__VDD_8 0.603529
R_x3_PM_AND2_X2__VDD_r8 x3_PM_AND2_X2__VDD_17 x3_PM_AND2_X2__VDD_7 0.0731438
R_x3_PM_AND2_X2__VDD_r9 VDD x3_PM_AND2_X2__VDD_7 0.0894118
R_x3_PM_AND2_X2__VDD_r10 x3_PM_AND2_X2__VDD_8 x3_PM_AND2_X2__VDD_3 0.264221
R_x3_PM_AND2_X2__VDD_r11 N3_VDD_M0_s x3_PM_AND2_X2__VDD_3 0.420714
C_x3_PM_AND2_X2__3_c0 VSS x3_PM_AND2_X2__3_33 1.13133e-17
C_x3_PM_AND2_X2__3_c1 VSS x3_PM_AND2_X2__3_30 1.00152e-17
C_x3_PM_AND2_X2__3_c2 VSS x3_PM_AND2_X2__3_29 9.34287e-17
C_x3_PM_AND2_X2__3_c3 VSS x3_PM_AND2_X2__3_26 1.87365e-17
C_x3_PM_AND2_X2__3_c4 VSS x3_PM_AND2_X2__3_22 8.60574e-18
C_x3_PM_AND2_X2__3_c5 VSS x3_PM_AND2_X2__3_21 4.03179e-17
C_x3_PM_AND2_X2__3_c6 VSS N3_3_M0_d 3.31237e-17
C_x3_PM_AND2_X2__3_c7 VSS x3_PM_AND2_X2__3_16 5.73522e-18
C_x3_PM_AND2_X2__3_c8 VSS x3_PM_AND2_X2__3_15 6.02033e-17
C_x3_PM_AND2_X2__3_c9 VSS N3_3_M3_s 2.55776e-17
C_x3_PM_AND2_X2__3_c10 VSS N3_3_M2_g 9.71074e-17
C_x3_PM_AND2_X2__3_c11 VSS N3_3_M5_g 3.53623e-17
R_x3_PM_AND2_X2__3_r12 x3_PM_AND2_X2__3_33 x3_PM_AND2_X2__3_31 3.38
R_x3_PM_AND2_X2__3_r13 x3_PM_AND2_X2__3_29 x3_PM_AND2_X2__3_30 2.93143
R_x3_PM_AND2_X2__3_r14 x3_PM_AND2_X2__3_31 x3_PM_AND2_X2__3_26 25.0012
R_x3_PM_AND2_X2__3_r15 x3_PM_AND2_X2__3_30 x3_PM_AND2_X2__3_24 0.232321
R_x3_PM_AND2_X2__3_r16 x3_PM_AND2_X2__3_26 x3_PM_AND2_X2__3_24 0.0542857
R_x3_PM_AND2_X2__3_r17 x3_PM_AND2_X2__3_26 x3_PM_AND2_X2__3_23 0.22619
R_x3_PM_AND2_X2__3_r18 x3_PM_AND2_X2__3_29 x3_PM_AND2_X2__3_21 0.212317
R_x3_PM_AND2_X2__3_r19 x3_PM_AND2_X2__3_22 x3_PM_AND2_X2__3_21 0.76
R_x3_PM_AND2_X2__3_r20 x3_PM_AND2_X2__3_22 x3_PM_AND2_X2__3_17 0.212317
R_x3_PM_AND2_X2__3_r21 N3_3_M0_d x3_PM_AND2_X2__3_17 0.393571
R_x3_PM_AND2_X2__3_r22 x3_PM_AND2_X2__3_23 x3_PM_AND2_X2__3_15 0.223553
R_x3_PM_AND2_X2__3_r23 x3_PM_AND2_X2__3_16 x3_PM_AND2_X2__3_15 1.79143
R_x3_PM_AND2_X2__3_r24 x3_PM_AND2_X2__3_16 x3_PM_AND2_X2__3_11 0.212317
R_x3_PM_AND2_X2__3_r25 N3_3_M3_s x3_PM_AND2_X2__3_11 0.420714
R_x3_PM_AND2_X2__3_r26 x3_PM_AND2_X2__3_33 x3_PM_AND2_X2__3_5 1.95
R_x3_PM_AND2_X2__3_r27 N3_3_M2_g x3_PM_AND2_X2__3_5 105.3
R_x3_PM_AND2_X2__3_r28 x3_PM_AND2_X2__3_33 x3_PM_AND2_X2__3_VSS 1.95
R_x3_PM_AND2_X2__3_r29 N3_3_M5_g x3_PM_AND2_X2__3_VSS 27.3
C_x3_PM_AND2_X2__Zalp1_c0 VSS x3_PM_AND2_X2__Zalp1_13 7.02743e-18
C_x3_PM_AND2_X2__Zalp1_c1 VSS Zalp1 1.56682e-17
C_x3_PM_AND2_X2__Zalp1_c2 VSS N3_Zalp1_M0_g 6.18939e-17
C_x3_PM_AND2_X2__Zalp1_c3 VSS N3_Zalp1_M3_g 5.49708e-17
R_x3_PM_AND2_X2__Zalp1_r4 x3_PM_AND2_X2__Zalp1_16 x3_PM_AND2_X2__Zalp1_13 4.74714
R_x3_PM_AND2_X2__Zalp1_r5 x3_PM_AND2_X2__Zalp1_15 x3_PM_AND2_X2__Zalp1_13 4.74714
R_x3_PM_AND2_X2__Zalp1_r6 x3_PM_AND2_X2__Zalp1_13 x3_PM_AND2_X2__Zalp1_11 25.0012
R_x3_PM_AND2_X2__Zalp1_r7 x3_PM_AND2_X2__Zalp1_11 Zalp1 0.158563
R_x3_PM_AND2_X2__Zalp1_r8 N3_Zalp1_M0_g x3_PM_AND2_X2__Zalp1_16 83.85
R_x3_PM_AND2_X2__Zalp1_r9 N3_Zalp1_M3_g x3_PM_AND2_X2__Zalp1_15 63.18
C_x3_PM_AND2_X2__Zalp2_c0 VSS x3_PM_AND2_X2__Zalp2_14 8.64377e-18
C_x3_PM_AND2_X2__Zalp2_c1 VSS x3_PM_AND2_X2__Zalp2_12 4.37781e-17
C_x3_PM_AND2_X2__Zalp2_c2 VSS N3_Zalp2_M1_g 5.57959e-17
C_x3_PM_AND2_X2__Zalp2_c3 VSS N3_Zalp2_M4_g 7.00537e-17
R_x3_PM_AND2_X2__Zalp2_r4 x3_PM_AND2_X2__Zalp2_18 x3_PM_AND2_X2__Zalp2_14 4.7687
R_x3_PM_AND2_X2__Zalp2_r5 x3_PM_AND2_X2__Zalp2_17 x3_PM_AND2_X2__Zalp2_14 4.7687
R_x3_PM_AND2_X2__Zalp2_r6 x3_PM_AND2_X2__Zalp2_14 x3_PM_AND2_X2__Zalp2_12 25.0012
R_x3_PM_AND2_X2__Zalp2_r7 x3_PM_AND2_X2__Zalp2_12 Zalp2 0.169643
R_x3_PM_AND2_X2__Zalp2_r8 N3_Zalp2_M1_g x3_PM_AND2_X2__Zalp2_18 62.01
R_x3_PM_AND2_X2__Zalp2_r9 N3_Zalp2_M4_g x3_PM_AND2_X2__Zalp2_17 85.02
C_x3_PM_AND2_X2__ZN3_c0 VSS N3_ZN3_M5_d 2.60988e-17
C_x3_PM_AND2_X2__ZN3_c1 VSS ZN 7.63258e-17
C_x3_PM_AND2_X2__ZN3_c2 VSS N3_ZN3_M2_d 5.16564e-17
C_x3_PM_AND2_X2__ZN3_c3 VSS x3_PM_AND2_X2__ZN3_3 6.61381e-18
R_x3_PM_AND2_X2__ZN3_r4 ZN x3_PM_AND2_X2__ZN3_8 1.87286
R_x3_PM_AND2_X2__ZN3_r5 x3_PM_AND2_X2__ZN3_7 N3_ZN3_M5_d 0.30478
R_x3_PM_AND2_X2__ZN3_r6 ZN x3_PM_AND2_X2__ZN3_7 1.60143
R_x3_PM_AND2_X2__ZN3_r7 x3_PM_AND2_X2__ZN3_8 x3_PM_AND2_X2__ZN3_3 0.20978
R_x3_PM_AND2_X2__ZN3_r8 N3_ZN3_M2_d x3_PM_AND2_X2__ZN3_3 0.686111
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
