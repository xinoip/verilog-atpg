.SUBCKT buf1 A VDD VSS Z 
M_M2 N_VDD_M0_d N_A_M0_g N_3_M0_s VDD PMOS_VTL L=0.050U W=0.135000U AS=0.014175P AD=0.028350P PS=0.480000U PD=0.820000U
M_M3 N_Z_M1_d N_3_M1_g N_VDD_M0_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 N_VSS_M2_d N_A_M2_g N_3_M2_s VSS NMOS_VTL L=0.050U W=0.090000U AS=0.009450P AD=0.018900P PS=0.390000U PD=0.640000U
M_M1 N_Z_M3_d N_3_M3_g N_VSS_M2_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_BUF_X2__VSS_c0 VSS VSS 1.0786e-16
R_x_PM_BUF_X2__VSS_r1 N_VSS_M2_d VSS 0.637857
C_x_PM_BUF_X2__VDD_c0 VSS VDD 8.03115e-17
C_x_PM_BUF_X2__VDD_c1 VSS N_VDD_M0_d 3.78724e-17
R_x_PM_BUF_X2__VDD_r2 VDD x_PM_BUF_X2__VDD_4 0.145286
R_x_PM_BUF_X2__VDD_r3 N_VDD_M0_d x_PM_BUF_X2__VDD_4 0.420714
C_x_PM_BUF_X2__3_c0 VSS x_PM_BUF_X2__3_31 9.87551e-18
C_x_PM_BUF_X2__3_c1 VSS x_PM_BUF_X2__3_25 4.34052e-17
C_x_PM_BUF_X2__3_c2 VSS x_PM_BUF_X2__3_24 9.58887e-17
C_x_PM_BUF_X2__3_c3 VSS x_PM_BUF_X2__3_22 4.39826e-18
C_x_PM_BUF_X2__3_c4 VSS x_PM_BUF_X2__3_21 4.41595e-17
C_x_PM_BUF_X2__3_c5 VSS x_PM_BUF_X2__3_20 1.51022e-17
C_x_PM_BUF_X2__3_c6 VSS x_PM_BUF_X2__3_19 2.89567e-17
C_x_PM_BUF_X2__3_c7 VSS N_3_M0_s 2.73356e-17
C_x_PM_BUF_X2__3_c8 VSS N_3_M2_s 3.67549e-17
C_x_PM_BUF_X2__3_c9 VSS N_3_M1_g 8.56064e-17
C_x_PM_BUF_X2__3_c10 VSS N_3_M3_g 4.79448e-17
R_x_PM_BUF_X2__3_r11 x_PM_BUF_X2__3_33 x_PM_BUF_X2__3_31 4.74714
R_x_PM_BUF_X2__3_r12 x_PM_BUF_X2__3_30 x_PM_BUF_X2__3_28 0.297071
R_x_PM_BUF_X2__3_r13 x_PM_BUF_X2__3_31 x_PM_BUF_X2__3_28 25.0012
R_x_PM_BUF_X2__3_r14 x_PM_BUF_X2__3_28 x_PM_BUF_X2__3_25 0.13
R_x_PM_BUF_X2__3_r15 x_PM_BUF_X2__3_24 x_PM_BUF_X2__3_30 2.57857
R_x_PM_BUF_X2__3_r16 x_PM_BUF_X2__3_24 x_PM_BUF_X2__3_21 0.212317
R_x_PM_BUF_X2__3_r17 x_PM_BUF_X2__3_22 x_PM_BUF_X2__3_21 0.895714
R_x_PM_BUF_X2__3_r18 x_PM_BUF_X2__3_25 x_PM_BUF_X2__3_19 0.095
R_x_PM_BUF_X2__3_r19 x_PM_BUF_X2__3_20 x_PM_BUF_X2__3_19 0.895714
R_x_PM_BUF_X2__3_r20 x_PM_BUF_X2__3_22 x_PM_BUF_X2__3_15 0.212317
R_x_PM_BUF_X2__3_r21 N_3_M0_s x_PM_BUF_X2__3_15 0.393571
R_x_PM_BUF_X2__3_r22 x_PM_BUF_X2__3_20 x_PM_BUF_X2__3_11 0.212317
R_x_PM_BUF_X2__3_r23 N_3_M2_s x_PM_BUF_X2__3_11 1.045
R_x_PM_BUF_X2__3_r24 N_3_M1_g x_PM_BUF_X2__3_33 95.16
R_x_PM_BUF_X2__3_r25 x_PM_BUF_X2__3_VSS x_PM_BUF_X2__3_31 4.74714
R_x_PM_BUF_X2__3_r26 N_3_M3_g x_PM_BUF_X2__3_VSS 42.9
C_x_PM_BUF_X2__A_c0 VSS x_PM_BUF_X2__A_14 7.38755e-18
C_x_PM_BUF_X2__A_c1 VSS x_PM_BUF_X2__A_12 6.51234e-17
C_x_PM_BUF_X2__A_c2 VSS N_A_M0_g 6.60639e-17
C_x_PM_BUF_X2__A_c3 VSS N_A_M2_g 5.42189e-17
R_x_PM_BUF_X2__A_r4 x_PM_BUF_X2__A_18 x_PM_BUF_X2__A_14 4.7687
R_x_PM_BUF_X2__A_r5 x_PM_BUF_X2__A_17 x_PM_BUF_X2__A_14 4.7687
R_x_PM_BUF_X2__A_r6 x_PM_BUF_X2__A_14 x_PM_BUF_X2__A_12 25.0012
R_x_PM_BUF_X2__A_r7 x_PM_BUF_X2__A_12 A 0.2375
R_x_PM_BUF_X2__A_r8 N_A_M0_g x_PM_BUF_X2__A_18 84.63
R_x_PM_BUF_X2__A_r9 N_A_M2_g x_PM_BUF_X2__A_17 56.94
C_x_PM_BUF_X2__Z_c0 VSS N_Z_M3_d 3.4635e-17
C_x_PM_BUF_X2__Z_c1 VSS Z 9.23569e-17
C_x_PM_BUF_X2__Z_c2 VSS N_Z_M1_d 5.59233e-17
C_x_PM_BUF_X2__Z_c3 VSS x_PM_BUF_X2__Z_3 8.95839e-18
R_x_PM_BUF_X2__Z_r4 Z x_PM_BUF_X2__Z_8 1.87286
R_x_PM_BUF_X2__Z_r5 x_PM_BUF_X2__Z_7 N_Z_M3_d 0.30478
R_x_PM_BUF_X2__Z_r6 Z x_PM_BUF_X2__Z_7 1.79143
R_x_PM_BUF_X2__Z_r7 x_PM_BUF_X2__Z_8 x_PM_BUF_X2__Z_3 0.20978
R_x_PM_BUF_X2__Z_r8 N_Z_M1_d x_PM_BUF_X2__Z_3 0.686111
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
