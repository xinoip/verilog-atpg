.SUBCKT nand3 A1 A2 A3 VDD VSS ZN 
M_M3 N_ZN_M0_d N_A3_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.037800P PS=0.750000U PD=0.820000U
M_M4 N_VDD_M1_d N_A2_M1_g N_ZN_M0_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.037800P PS=0.820000U PD=0.820000U
M_M5 N_ZN_M2_d N_A1_M2_g N_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 7 N_A3_M3_g N_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.340000U AS=0.035700P AD=0.047600P PS=0.890000U PD=0.960000U
M_M1 8 N_A2_M4_g 7 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.047600P PS=0.960000U PD=0.960000U
M_M2 N_ZN_M5_d N_A1_M5_g 8 VSS NMOS_VTL W=0.340000U AS=0.047600P AD=0.035700P PS=0.960000U PD=0.890000U
C_x_PM_NAND3_X2__VSS_c0 VSS VSS 7.02872e-17
C_x_PM_NAND3_X2__VSS_c1 VSS x_PM_NAND3_X2__VSS_6 1.05487e-17
C_x_PM_NAND3_X2__VSS_c2 VSS N_VSS_M3_s 1.8134e-17
R_x_PM_NAND3_X2__VSS_r3 VSS x_PM_NAND3_X2__VSS_6 0.603529
R_x_PM_NAND3_X2__VSS_r4 x_PM_NAND3_X2__VSS_6 x_PM_NAND3_X2__VSS_2 0.264221
R_x_PM_NAND3_X2__VSS_r5 N_VSS_M3_s x_PM_NAND3_X2__VSS_2 0.230714
C_x_PM_NAND3_X2__VDD_c0 VSS N_VDD_M1_d 6.12848e-17
C_x_PM_NAND3_X2__VDD_c1 VSS x_PM_NAND3_X2__VDD_7 3.00804e-17
C_x_PM_NAND3_X2__VDD_c2 VSS N_VDD_M0_s 2.5125e-17
C_x_PM_NAND3_X2__VDD_c3 VSS x_PM_NAND3_X2__VDD_3 1.06055e-17
R_x_PM_NAND3_X2__VDD_r4 VDD x_PM_NAND3_X2__VDD_8 0.195294
R_x_PM_NAND3_X2__VDD_r5 x_PM_NAND3_X2__VDD_7 N_VDD_M1_d 0.140674
R_x_PM_NAND3_X2__VDD_r6 x_PM_NAND3_X2__VDD_8 x_PM_NAND3_X2__VDD_7 0.614706
R_x_PM_NAND3_X2__VDD_r7 VDD x_PM_NAND3_X2__VDD_3 0.0689273
R_x_PM_NAND3_X2__VDD_r8 N_VDD_M0_s x_PM_NAND3_X2__VDD_3 0.230714
C_x_PM_NAND3_X2__A3_c0 VSS x_PM_NAND3_X2__A3_14 6.68331e-18
C_x_PM_NAND3_X2__A3_c1 VSS x_PM_NAND3_X2__A3_12 3.18495e-17
C_x_PM_NAND3_X2__A3_c2 VSS N_A3_M0_g 7.81987e-17
C_x_PM_NAND3_X2__A3_c3 VSS N_A3_M3_g 4.14029e-17
R_x_PM_NAND3_X2__A3_r4 x_PM_NAND3_X2__A3_18 x_PM_NAND3_X2__A3_14 4.7687
R_x_PM_NAND3_X2__A3_r5 x_PM_NAND3_X2__A3_17 x_PM_NAND3_X2__A3_14 4.7687
R_x_PM_NAND3_X2__A3_r6 x_PM_NAND3_X2__A3_14 x_PM_NAND3_X2__A3_12 25.0012
R_x_PM_NAND3_X2__A3_r7 x_PM_NAND3_X2__A3_12 A3 0.0781486
R_x_PM_NAND3_X2__A3_r8 N_A3_M0_g x_PM_NAND3_X2__A3_18 95.94
R_x_PM_NAND3_X2__A3_r9 N_A3_M3_g x_PM_NAND3_X2__A3_17 35.1
C_x_PM_NAND3_X2__ZN_c0 VSS N_ZN_M5_d 1.32739e-16
C_x_PM_NAND3_X2__ZN_c1 VSS x_PM_NAND3_X2__ZN_8 1.01878e-17
C_x_PM_NAND3_X2__ZN_c2 VSS x_PM_NAND3_X2__ZN_4 7.15422e-17
R_x_PM_NAND3_X2__ZN_r3 ZN N_ZN_M5_d 1.59389
R_x_PM_NAND3_X2__ZN_r4 N_ZN_M2_d x_PM_NAND3_X2__ZN_8 0.0406238
R_x_PM_NAND3_X2__ZN_r5 ZN x_PM_NAND3_X2__ZN_8 1.28778
R_x_PM_NAND3_X2__ZN_r6 N_ZN_M2_d x_PM_NAND3_X2__ZN_4 0.176037
R_x_PM_NAND3_X2__ZN_r7 N_ZN_M0_d x_PM_NAND3_X2__ZN_4 1.85929
C_x_PM_NAND3_X2__A2_c0 VSS x_PM_NAND3_X2__A2_14 8.63262e-18
C_x_PM_NAND3_X2__A2_c1 VSS x_PM_NAND3_X2__A2_12 3.91329e-17
C_x_PM_NAND3_X2__A2_c2 VSS N_A2_M1_g 4.24405e-17
C_x_PM_NAND3_X2__A2_c3 VSS N_A2_M4_g 8.48173e-17
R_x_PM_NAND3_X2__A2_r4 x_PM_NAND3_X2__A2_18 x_PM_NAND3_X2__A2_14 4.7687
R_x_PM_NAND3_X2__A2_r5 x_PM_NAND3_X2__A2_17 x_PM_NAND3_X2__A2_14 4.7687
R_x_PM_NAND3_X2__A2_r6 x_PM_NAND3_X2__A2_14 x_PM_NAND3_X2__A2_12 25.0012
R_x_PM_NAND3_X2__A2_r7 x_PM_NAND3_X2__A2_12 A2 0.169643
R_x_PM_NAND3_X2__A2_r8 N_A2_M1_g x_PM_NAND3_X2__A2_18 29.64
R_x_PM_NAND3_X2__A2_r9 N_A2_M4_g x_PM_NAND3_X2__A2_17 101.4
C_x_PM_NAND3_X2__A1_c0 VSS x_PM_NAND3_X2__A1_18 1.22048e-17
C_x_PM_NAND3_X2__A1_c1 VSS x_PM_NAND3_X2__A1_12 7.61168e-17
C_x_PM_NAND3_X2__A1_c2 VSS N_A1_M2_g 8.98944e-17
C_x_PM_NAND3_X2__A1_c3 VSS N_A1_M5_g 4.86035e-17
R_x_PM_NAND3_X2__A1_r4 x_PM_NAND3_X2__A1_18 x_PM_NAND3_X2__A1_14 3.9
R_x_PM_NAND3_X2__A1_r5 x_PM_NAND3_X2__A1_14 x_PM_NAND3_X2__A1_12 25.0012
R_x_PM_NAND3_X2__A1_r6 x_PM_NAND3_X2__A1_12 A1 0.0459677
R_x_PM_NAND3_X2__A1_r7 x_PM_NAND3_X2__A1_18 x_PM_NAND3_X2__A1_5 1.95
R_x_PM_NAND3_X2__A1_r8 N_A1_M2_g x_PM_NAND3_X2__A1_5 95.94
R_x_PM_NAND3_X2__A1_r9 x_PM_NAND3_X2__A1_18 x_PM_NAND3_X2__A1_VSS 1.95
R_x_PM_NAND3_X2__A1_r10 N_A1_M5_g x_PM_NAND3_X2__A1_VSS 35.1
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
