.SUBCKT nor3 A1 A2 A3 VDD VSS ZN 
M_M3 7 N_A3_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.520000U AS=0.054600P AD=0.072800P PS=1.250000U PD=1.320000U
M_M4 8 N_A2_M1_g 7 VDD PMOS_VTL L=0.050U W=0.520000U AS=0.072800P AD=0.072800P PS=1.320000U PD=1.320000U
M_M5 N_ZN_M2_d N_A1_M2_g 8 VDD PMOS_VTL L=0.050U W=0.520000U AS=0.072800P AD=0.054600P PS=1.320000U PD=1.250000U
M_M0 N_ZN_M3_d N_A3_M3_g N_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M_M1 N_VSS_M4_d N_A2_M4_g N_ZN_M3_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M_M2 N_ZN_M5_d N_A1_M5_g N_VSS_M4_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_NOR3_X2__VSS_c0 VSS x_PM_NOR3_X2__VSS_17 4.46075e-17
C_x_PM_NOR3_X2__VSS_c1 VSS N_VSS_M4_d 2.78358e-17
C_x_PM_NOR3_X2__VSS_c2 VSS x_PM_NOR3_X2__VSS_8 1.05487e-17
C_x_PM_NOR3_X2__VSS_c3 VSS x_PM_NOR3_X2__VSS_7 3.86305e-17
C_x_PM_NOR3_X2__VSS_c4 VSS N_VSS_M3_s 9.87304e-18
R_x_PM_NOR3_X2__VSS_r5 x_PM_NOR3_X2__VSS_17 x_PM_NOR3_X2__VSS_11 0.145286
R_x_PM_NOR3_X2__VSS_r6 N_VSS_M4_d x_PM_NOR3_X2__VSS_11 0.230714
R_x_PM_NOR3_X2__VSS_r7 VSS x_PM_NOR3_X2__VSS_8 0.603529
R_x_PM_NOR3_X2__VSS_r8 x_PM_NOR3_X2__VSS_17 x_PM_NOR3_X2__VSS_7 0.0731438
R_x_PM_NOR3_X2__VSS_r9 VSS x_PM_NOR3_X2__VSS_7 0.0782353
R_x_PM_NOR3_X2__VSS_r10 x_PM_NOR3_X2__VSS_8 x_PM_NOR3_X2__VSS_3 0.264221
R_x_PM_NOR3_X2__VSS_r11 N_VSS_M3_s x_PM_NOR3_X2__VSS_3 0.230714
C_x_PM_NOR3_X2__VDD_c0 VSS VDD 5.9596e-17
C_x_PM_NOR3_X2__VDD_c1 VSS N_VDD_M0_s 2.58417e-17
C_x_PM_NOR3_X2__VDD_c2 VSS x_PM_NOR3_X2__VDD_2 1.06055e-17
R_x_PM_NOR3_X2__VDD_r3 VDD x_PM_NOR3_X2__VDD_2 0.0689273
R_x_PM_NOR3_X2__VDD_r4 N_VDD_M0_s x_PM_NOR3_X2__VDD_2 0.230714
C_x_PM_NOR3_X2__A3_c0 VSS x_PM_NOR3_X2__A3_11 7.14715e-18
C_x_PM_NOR3_X2__A3_c1 VSS x_PM_NOR3_X2__A3_9 5.04542e-17
C_x_PM_NOR3_X2__A3_c2 VSS N_A3_M0_g 6.20936e-17
C_x_PM_NOR3_X2__A3_c3 VSS N_A3_M3_g 5.91756e-17
R_x_PM_NOR3_X2__A3_r4 x_PM_NOR3_X2__A3_18 x_PM_NOR3_X2__A3_11 4.74714
R_x_PM_NOR3_X2__A3_r5 x_PM_NOR3_X2__A3_17 x_PM_NOR3_X2__A3_11 4.74714
R_x_PM_NOR3_X2__A3_r6 x_PM_NOR3_X2__A3_11 x_PM_NOR3_X2__A3_9 25.0012
R_x_PM_NOR3_X2__A3_r7 A3 x_PM_NOR3_X2__A3_9 0.2204
R_x_PM_NOR3_X2__A3_r8 N_A3_M0_g x_PM_NOR3_X2__A3_18 49.14
R_x_PM_NOR3_X2__A3_r9 N_A3_M3_g x_PM_NOR3_X2__A3_17 74.88
C_x_PM_NOR3_X2__ZN_c0 VSS x_PM_NOR3_X2__ZN_22 2.56413e-18
C_x_PM_NOR3_X2__ZN_c1 VSS ZN 5.06951e-17
C_x_PM_NOR3_X2__ZN_c2 VSS N_ZN_M2_d 2.75881e-17
C_x_PM_NOR3_X2__ZN_c3 VSS x_PM_NOR3_X2__ZN_14 6.25994e-18
C_x_PM_NOR3_X2__ZN_c4 VSS N_ZN_M5_d 2.52851e-17
C_x_PM_NOR3_X2__ZN_c5 VSS x_PM_NOR3_X2__ZN_9 8.16416e-18
C_x_PM_NOR3_X2__ZN_c6 VSS x_PM_NOR3_X2__ZN_8 4.12951e-17
C_x_PM_NOR3_X2__ZN_c7 VSS N_ZN_M3_d 2.15312e-17
R_x_PM_NOR3_X2__ZN_r8 ZN x_PM_NOR3_X2__ZN_19 1.46571
R_x_PM_NOR3_X2__ZN_r9 x_PM_NOR3_X2__ZN_22 x_PM_NOR3_X2__ZN_18 0.143785
R_x_PM_NOR3_X2__ZN_r10 ZN x_PM_NOR3_X2__ZN_18 0.868571
R_x_PM_NOR3_X2__ZN_r11 x_PM_NOR3_X2__ZN_19 x_PM_NOR3_X2__ZN_14 0.20978
R_x_PM_NOR3_X2__ZN_r12 N_ZN_M2_d x_PM_NOR3_X2__ZN_14 0.686111
R_x_PM_NOR3_X2__ZN_r13 x_PM_NOR3_X2__ZN_22 x_PM_NOR3_X2__ZN_10 0.143785
R_x_PM_NOR3_X2__ZN_r14 N_ZN_M5_d x_PM_NOR3_X2__ZN_10 0.116111
R_x_PM_NOR3_X2__ZN_r15 x_PM_NOR3_X2__ZN_22 x_PM_NOR3_X2__ZN_8 0.0569232
R_x_PM_NOR3_X2__ZN_r16 x_PM_NOR3_X2__ZN_9 x_PM_NOR3_X2__ZN_8 1.65571
R_x_PM_NOR3_X2__ZN_r17 x_PM_NOR3_X2__ZN_9 x_PM_NOR3_X2__ZN_4 0.212317
R_x_PM_NOR3_X2__ZN_r18 N_ZN_M3_d x_PM_NOR3_X2__ZN_4 0.149286
C_x_PM_NOR3_X2__A2_c0 VSS x_PM_NOR3_X2__A2_11 8.98632e-18
C_x_PM_NOR3_X2__A2_c1 VSS x_PM_NOR3_X2__A2_9 8.53584e-17
C_x_PM_NOR3_X2__A2_c2 VSS N_A2_M1_g 6.12109e-17
C_x_PM_NOR3_X2__A2_c3 VSS N_A2_M4_g 6.60015e-17
R_x_PM_NOR3_X2__A2_r4 x_PM_NOR3_X2__A2_18 x_PM_NOR3_X2__A2_11 4.74714
R_x_PM_NOR3_X2__A2_r5 x_PM_NOR3_X2__A2_17 x_PM_NOR3_X2__A2_11 4.74714
R_x_PM_NOR3_X2__A2_r6 x_PM_NOR3_X2__A2_11 x_PM_NOR3_X2__A2_9 25.0012
R_x_PM_NOR3_X2__A2_r7 A2 x_PM_NOR3_X2__A2_9 0.2204
R_x_PM_NOR3_X2__A2_r8 N_A2_M1_g x_PM_NOR3_X2__A2_18 49.14
R_x_PM_NOR3_X2__A2_r9 N_A2_M4_g x_PM_NOR3_X2__A2_17 74.88
C_x_PM_NOR3_X2__A1_c0 VSS x_PM_NOR3_X2__A1_20 1.07269e-17
C_x_PM_NOR3_X2__A1_c1 VSS x_PM_NOR3_X2__A1_14 4.59258e-17
C_x_PM_NOR3_X2__A1_c2 VSS x_PM_NOR3_X2__A1_9 3.45973e-17
C_x_PM_NOR3_X2__A1_c3 VSS N_A1_M2_g 7.00434e-17
C_x_PM_NOR3_X2__A1_c4 VSS N_A1_M5_g 6.63408e-17
R_x_PM_NOR3_X2__A1_r5 x_PM_NOR3_X2__A1_20 x_PM_NOR3_X2__A1_16 2.34
R_x_PM_NOR3_X2__A1_r6 x_PM_NOR3_X2__A1_16 x_PM_NOR3_X2__A1_14 25.0012
R_x_PM_NOR3_X2__A1_r7 x_PM_NOR3_X2__A1_14 x_PM_NOR3_X2__A1_12 0.147778
R_x_PM_NOR3_X2__A1_r8 x_PM_NOR3_X2__A1_12 x_PM_NOR3_X2__A1_9 0.095
R_x_PM_NOR3_X2__A1_r9 A1 x_PM_NOR3_X2__A1_9 0.298571
R_x_PM_NOR3_X2__A1_r10 x_PM_NOR3_X2__A1_20 x_PM_NOR3_X2__A1_5 1.95
R_x_PM_NOR3_X2__A1_r11 N_A1_M2_g x_PM_NOR3_X2__A1_5 56.94
R_x_PM_NOR3_X2__A1_r12 x_PM_NOR3_X2__A1_20 x_PM_NOR3_X2__A1_VSS 1.95
R_x_PM_NOR3_X2__A1_r13 N_A1_M5_g x_PM_NOR3_X2__A1_VSS 67.08
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
