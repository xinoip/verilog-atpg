.SUBCKT or4 A1 A2 A3 A4 VDD VSS ZN 
M_M5 9 N_A1_M0_g N_3_M0_s VDD PMOS_VTL L=0.050U W=0.325000U AS=0.034125P AD=0.045500P PS=0.860000U PD=0.930000U
M_M6 10 N_A2_M1_g 9 VDD PMOS_VTL L=0.050U W=0.325000U AS=0.045500P AD=0.045500P PS=0.930000U PD=0.930000U
M_M7 11 N_A3_M2_g 10 VDD PMOS_VTL L=0.050U W=0.325000U AS=0.045500P AD=0.045500P PS=0.930000U PD=0.930000U
M_M8 N_VDD_M3_d N_A4_M3_g 11 VDD PMOS_VTL L=0.050U W=0.325000U AS=0.045500P AD=0.041650P PS=0.930000U PD=0.930000U
M_M9 N_ZN_M4_d N_3_M4_g N_VDD_M3_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.041650P AD=0.028350P PS=0.930000U PD=0.750000U
M_M0 N_3_M5_d N_A1_M5_g N_VSS_M5_s VSS NMOS_VTL L=0.050U W=0.090000U AS=0.009450P AD=0.012600P PS=0.390000U PD=0.460000U
M_M1 N_VSS_M6_d N_A2_M6_g N_3_M5_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.012600P PS=0.460000U PD=0.460000U
M_M2 N_3_M7_d N_A3_M7_g N_VSS_M6_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.012600P PS=0.460000U PD=0.460000U
M_M3 N_VSS_M8_d N_A4_M8_g N_3_M7_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.018900P PS=0.460000U PD=0.600000U
M_M4 N_ZN_M9_d N_3_M9_g N_VSS_M8_d VSS NMOS_VTL L=0.050U W=0.160000U AS=0.018900P AD=0.020000P PS=0.600000U PD=0.570000U
C_x_PM_OR4_X2__VSS_c0 VSS x_PM_OR4_X2__VSS_25 3.09849e-17
C_x_PM_OR4_X2__VSS_c1 VSS x_PM_OR4_X2__VSS_24 2.92048e-18
C_x_PM_OR4_X2__VSS_c2 VSS N_VSS_M8_d 3.12663e-17
C_x_PM_OR4_X2__VSS_c3 VSS x_PM_OR4_X2__VSS_14 3.18026e-17
C_x_PM_OR4_X2__VSS_c4 VSS N_VSS_M6_d 3.20111e-17
C_x_PM_OR4_X2__VSS_c5 VSS x_PM_OR4_X2__VSS_9 1.25763e-17
C_x_PM_OR4_X2__VSS_c6 VSS x_PM_OR4_X2__VSS_8 3.12295e-17
C_x_PM_OR4_X2__VSS_c7 VSS N_VSS_M5_s 2.60989e-17
R_x_PM_OR4_X2__VSS_r8 x_PM_OR4_X2__VSS_25 x_PM_OR4_X2__VSS_18 0.145286
R_x_PM_OR4_X2__VSS_r9 N_VSS_M8_d x_PM_OR4_X2__VSS_18 0.637857
R_x_PM_OR4_X2__VSS_r10 x_PM_OR4_X2__VSS_24 x_PM_OR4_X2__VSS_15 0.0731438
R_x_PM_OR4_X2__VSS_r11 VSS x_PM_OR4_X2__VSS_15 0.145294
R_x_PM_OR4_X2__VSS_r12 x_PM_OR4_X2__VSS_25 x_PM_OR4_X2__VSS_14 0.0731438
R_x_PM_OR4_X2__VSS_r13 VSS x_PM_OR4_X2__VSS_14 0.547647
R_x_PM_OR4_X2__VSS_r14 x_PM_OR4_X2__VSS_24 x_PM_OR4_X2__VSS_10 0.145286
R_x_PM_OR4_X2__VSS_r15 N_VSS_M6_d x_PM_OR4_X2__VSS_10 0.637857
R_x_PM_OR4_X2__VSS_r16 x_PM_OR4_X2__VSS_24 x_PM_OR4_X2__VSS_8 0.0731438
R_x_PM_OR4_X2__VSS_r17 x_PM_OR4_X2__VSS_9 x_PM_OR4_X2__VSS_8 0.681765
R_x_PM_OR4_X2__VSS_r18 x_PM_OR4_X2__VSS_9 x_PM_OR4_X2__VSS_4 0.264221
R_x_PM_OR4_X2__VSS_r19 N_VSS_M5_s x_PM_OR4_X2__VSS_4 0.637857
C_x_PM_OR4_X2__VDD_c0 VSS x_PM_OR4_X2__VDD_12 2.87042e-17
C_x_PM_OR4_X2__VDD_c1 VSS N_VDD_M3_d 3.86698e-17
C_x_PM_OR4_X2__VDD_c2 VSS x_PM_OR4_X2__VDD_2 8.27814e-17
R_x_PM_OR4_X2__VDD_r3 x_PM_OR4_X2__VDD_12 x_PM_OR4_X2__VDD_6 0.145286
R_x_PM_OR4_X2__VDD_r4 N_VDD_M3_d x_PM_OR4_X2__VDD_6 0.529286
R_x_PM_OR4_X2__VDD_r5 x_PM_OR4_X2__VDD_12 x_PM_OR4_X2__VDD_2 0.0731438
R_x_PM_OR4_X2__VDD_r6 VDD x_PM_OR4_X2__VDD_2 0.910882
C_x_PM_OR4_X2__3_c0 VSS x_PM_OR4_X2__3_39 1.50137e-17
C_x_PM_OR4_X2__3_c1 VSS x_PM_OR4_X2__3_34 5.66088e-17
C_x_PM_OR4_X2__3_c2 VSS x_PM_OR4_X2__3_31 7.64543e-18
C_x_PM_OR4_X2__3_c3 VSS N_3_M7_d 4.36971e-17
C_x_PM_OR4_X2__3_c4 VSS x_PM_OR4_X2__3_24 3.90305e-17
C_x_PM_OR4_X2__3_c5 VSS N_3_M5_d 4.58822e-17
C_x_PM_OR4_X2__3_c6 VSS x_PM_OR4_X2__3_19 1.0509e-17
C_x_PM_OR4_X2__3_c7 VSS x_PM_OR4_X2__3_18 1.72682e-17
C_x_PM_OR4_X2__3_c8 VSS N_3_M0_s 3.58537e-17
C_x_PM_OR4_X2__3_c9 VSS x_PM_OR4_X2__3_14 4.30213e-18
C_x_PM_OR4_X2__3_c10 VSS x_PM_OR4_X2__3_13 5.51576e-17
C_x_PM_OR4_X2__3_c11 VSS N_3_M4_g 9.51623e-17
C_x_PM_OR4_X2__3_c12 VSS N_3_M9_g 3.01638e-17
R_x_PM_OR4_X2__3_r13 x_PM_OR4_X2__3_39 x_PM_OR4_X2__3_37 5.46
R_x_PM_OR4_X2__3_r14 x_PM_OR4_X2__3_37 x_PM_OR4_X2__3_34 25.0012
R_x_PM_OR4_X2__3_r15 x_PM_OR4_X2__3_34 x_PM_OR4_X2__3_32 1.28929
R_x_PM_OR4_X2__3_r16 x_PM_OR4_X2__3_32 x_PM_OR4_X2__3_26 0.095
R_x_PM_OR4_X2__3_r17 N_3_M7_d x_PM_OR4_X2__3_26 0.855
R_x_PM_OR4_X2__3_r18 x_PM_OR4_X2__3_31 x_PM_OR4_X2__3_25 0.160909
R_x_PM_OR4_X2__3_r19 x_PM_OR4_X2__3_32 x_PM_OR4_X2__3_24 0.19
R_x_PM_OR4_X2__3_r20 x_PM_OR4_X2__3_25 x_PM_OR4_X2__3_24 1.68286
R_x_PM_OR4_X2__3_r21 x_PM_OR4_X2__3_31 x_PM_OR4_X2__3_20 0.0418175
R_x_PM_OR4_X2__3_r22 N_3_M5_d x_PM_OR4_X2__3_20 0.855
R_x_PM_OR4_X2__3_r23 x_PM_OR4_X2__3_31 x_PM_OR4_X2__3_18 0.160909
R_x_PM_OR4_X2__3_r24 x_PM_OR4_X2__3_19 x_PM_OR4_X2__3_18 0.76
R_x_PM_OR4_X2__3_r25 N_3_M0_s x_PM_OR4_X2__3_14 0.64
R_x_PM_OR4_X2__3_r26 x_PM_OR4_X2__3_13 x_PM_OR4_X2__3_14 0.217071
R_x_PM_OR4_X2__3_r27 x_PM_OR4_X2__3_19 x_PM_OR4_X2__3_12 0.212317
R_x_PM_OR4_X2__3_r28 x_PM_OR4_X2__3_13 x_PM_OR4_X2__3_12 2.76857
R_x_PM_OR4_X2__3_r29 x_PM_OR4_X2__3_39 x_PM_OR4_X2__3_5 1.95
R_x_PM_OR4_X2__3_r30 N_3_M4_g x_PM_OR4_X2__3_5 104.52
R_x_PM_OR4_X2__3_r31 x_PM_OR4_X2__3_39 x_PM_OR4_X2__3_VSS 1.95
R_x_PM_OR4_X2__3_r32 N_3_M9_g x_PM_OR4_X2__3_VSS 20.28
C_x_PM_OR4_X2__A1_c0 VSS A1 7.09523e-17
C_x_PM_OR4_X2__A1_c1 VSS x_PM_OR4_X2__A1_11 9.93232e-18
C_x_PM_OR4_X2__A1_c2 VSS N_A1_M0_g 7.76163e-17
C_x_PM_OR4_X2__A1_c3 VSS N_A1_M5_g 5.54373e-17
R_x_PM_OR4_X2__A1_r4 x_PM_OR4_X2__A1_18 x_PM_OR4_X2__A1_11 4.7687
R_x_PM_OR4_X2__A1_r5 x_PM_OR4_X2__A1_17 x_PM_OR4_X2__A1_11 4.7687
R_x_PM_OR4_X2__A1_r6 x_PM_OR4_X2__A1_11 x_PM_OR4_X2__A1_9 25.0012
R_x_PM_OR4_X2__A1_r7 A1 x_PM_OR4_X2__A1_9 0.223929
R_x_PM_OR4_X2__A1_r8 N_A1_M0_g x_PM_OR4_X2__A1_18 75.27
R_x_PM_OR4_X2__A1_r9 N_A1_M5_g x_PM_OR4_X2__A1_17 59.28
C_x_PM_OR4_X2__A2_c0 VSS A2 6.65609e-17
C_x_PM_OR4_X2__A2_c1 VSS x_PM_OR4_X2__A2_11 1.12437e-17
C_x_PM_OR4_X2__A2_c2 VSS N_A2_M1_g 6.83316e-17
C_x_PM_OR4_X2__A2_c3 VSS N_A2_M6_g 5.1084e-17
R_x_PM_OR4_X2__A2_r4 x_PM_OR4_X2__A2_11 x_PM_OR4_X2__A2_16 3.9
R_x_PM_OR4_X2__A2_r5 x_PM_OR4_X2__A2_11 x_PM_OR4_X2__A2_9 25.0012
R_x_PM_OR4_X2__A2_r6 A2 x_PM_OR4_X2__A2_9 0.156071
R_x_PM_OR4_X2__A2_r7 x_PM_OR4_X2__A2_16 x_PM_OR4_X2__A2_5 1.95
R_x_PM_OR4_X2__A2_r8 N_A2_M1_g x_PM_OR4_X2__A2_5 75.27
R_x_PM_OR4_X2__A2_r9 x_PM_OR4_X2__A2_16 x_PM_OR4_X2__A2_VSS 1.95
R_x_PM_OR4_X2__A2_r10 N_A2_M6_g x_PM_OR4_X2__A2_VSS 59.28
C_x_PM_OR4_X2__A3_c0 VSS A3 6.65126e-17
C_x_PM_OR4_X2__A3_c1 VSS x_PM_OR4_X2__A3_11 1.13495e-17
C_x_PM_OR4_X2__A3_c2 VSS N_A3_M2_g 6.82754e-17
C_x_PM_OR4_X2__A3_c3 VSS N_A3_M7_g 5.11699e-17
R_x_PM_OR4_X2__A3_r4 x_PM_OR4_X2__A3_11 x_PM_OR4_X2__A3_16 3.9
R_x_PM_OR4_X2__A3_r5 x_PM_OR4_X2__A3_11 x_PM_OR4_X2__A3_9 25.0012
R_x_PM_OR4_X2__A3_r6 A3 x_PM_OR4_X2__A3_9 0.156071
R_x_PM_OR4_X2__A3_r7 x_PM_OR4_X2__A3_16 x_PM_OR4_X2__A3_5 1.95
R_x_PM_OR4_X2__A3_r8 N_A3_M2_g x_PM_OR4_X2__A3_5 75.27
R_x_PM_OR4_X2__A3_r9 x_PM_OR4_X2__A3_16 x_PM_OR4_X2__A3_VSS 1.95
R_x_PM_OR4_X2__A3_r10 N_A3_M7_g x_PM_OR4_X2__A3_VSS 59.28
C_x_PM_OR4_X2__A4_c0 VSS A4 5.3212e-17
C_x_PM_OR4_X2__A4_c1 VSS x_PM_OR4_X2__A4_11 1.147e-17
C_x_PM_OR4_X2__A4_c2 VSS N_A4_M3_g 6.91639e-17
C_x_PM_OR4_X2__A4_c3 VSS N_A4_M8_g 5.25901e-17
R_x_PM_OR4_X2__A4_r4 x_PM_OR4_X2__A4_11 x_PM_OR4_X2__A4_16 3.9
R_x_PM_OR4_X2__A4_r5 x_PM_OR4_X2__A4_11 x_PM_OR4_X2__A4_9 25.0012
R_x_PM_OR4_X2__A4_r6 A4 x_PM_OR4_X2__A4_9 0.156071
R_x_PM_OR4_X2__A4_r7 x_PM_OR4_X2__A4_16 x_PM_OR4_X2__A4_5 1.95
R_x_PM_OR4_X2__A4_r8 N_A4_M3_g x_PM_OR4_X2__A4_5 75.27
R_x_PM_OR4_X2__A4_r9 x_PM_OR4_X2__A4_16 x_PM_OR4_X2__A4_VSS 1.95
R_x_PM_OR4_X2__A4_r10 N_A4_M8_g x_PM_OR4_X2__A4_VSS 59.28
C_x_PM_OR4_X2__ZN_c0 VSS N_ZN_M9_d 4.27646e-17
C_x_PM_OR4_X2__ZN_c1 VSS ZN 5.15232e-17
C_x_PM_OR4_X2__ZN_c2 VSS x_PM_OR4_X2__ZN_3 6.09228e-18
R_x_PM_OR4_X2__ZN_r3 N_ZN_M9_d x_PM_OR4_X2__ZN_13 1.47929
R_x_PM_OR4_X2__ZN_r4 N_ZN_M4_d ZN 1.65722
R_x_PM_OR4_X2__ZN_r5 x_PM_OR4_X2__ZN_13 x_PM_OR4_X2__ZN_3 0.20978
R_x_PM_OR4_X2__ZN_r6 ZN x_PM_OR4_X2__ZN_3 0.105556
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
