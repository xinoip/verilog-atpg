.SUBCKT or5 A1 A2 A3 A4 A5 VDD VSS ZN
********************************************NOR3_X2****************************************************
M_M3 7 N_A3_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.520000U AS=0.054600P AD=0.072800P PS=1.250000U PD=1.320000U
M_M4 8 N_A2_M1_g 7 VDD PMOS_VTL L=0.050U W=0.520000U AS=0.072800P AD=0.072800P PS=1.320000U PD=1.320000U
M_M5 N_Zalp1_M2_d N_A1_M2_g 8 VDD PMOS_VTL L=0.050U W=0.520000U AS=0.072800P AD=0.054600P PS=1.320000U PD=1.250000U
M_M0 N_Zalp1_M3_d N_A3_M3_g N_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M_M1 N_VSS_M4_d N_A2_M4_g N_Zalp1_M3_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M_M2 N_Zalp1_M5_d N_A1_M5_g N_VSS_M4_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_NOR3_X2__VSS_c0 VSS x_PM_NOR3_X2__VSS_17 4.46075e-17
C_x_PM_NOR3_X2__VSS_c1 VSS N_VSS_M4_d 2.78358e-17
C_x_PM_NOR3_X2__VSS_c2 VSS x_PM_NOR3_X2__VSS_8 1.05487e-17
C_x_PM_NOR3_X2__VSS_c3 VSS x_PM_NOR3_X2__VSS_7 3.86305e-17
C_x_PM_NOR3_X2__VSS_c4 VSS N_VSS_M3_s 9.87304e-18
R_x_PM_NOR3_X2__VSS_r5 x_PM_NOR3_X2__VSS_17 x_PM_NOR3_X2__VSS_11 0.145286
R_x_PM_NOR3_X2__VSS_r6 N_VSS_M4_d x_PM_NOR3_X2__VSS_11 0.230714
R_x_PM_NOR3_X2__VSS_r7 VSS x_PM_NOR3_X2__VSS_8 0.603529
R_x_PM_NOR3_X2__VSS_r8 x_PM_NOR3_X2__VSS_17 x_PM_NOR3_X2__VSS_7 0.0731438
R_x_PM_NOR3_X2__VSS_r9 VSS x_PM_NOR3_X2__VSS_7 0.0782353
R_x_PM_NOR3_X2__VSS_r10 x_PM_NOR3_X2__VSS_8 x_PM_NOR3_X2__VSS_3 0.264221
R_x_PM_NOR3_X2__VSS_r11 N_VSS_M3_s x_PM_NOR3_X2__VSS_3 0.230714
C_x_PM_NOR3_X2__VDD_c0 VSS VDD 5.9596e-17
C_x_PM_NOR3_X2__VDD_c1 VSS N_VDD_M0_s 2.58417e-17
C_x_PM_NOR3_X2__VDD_c2 VSS x_PM_NOR3_X2__VDD_2 1.06055e-17
R_x_PM_NOR3_X2__VDD_r3 VDD x_PM_NOR3_X2__VDD_2 0.0689273
R_x_PM_NOR3_X2__VDD_r4 N_VDD_M0_s x_PM_NOR3_X2__VDD_2 0.230714
C_x_PM_NOR3_X2__A3_c0 VSS x_PM_NOR3_X2__A3_11 7.14715e-18
C_x_PM_NOR3_X2__A3_c1 VSS x_PM_NOR3_X2__A3_9 5.04542e-17
C_x_PM_NOR3_X2__A3_c2 VSS N_A3_M0_g 6.20936e-17
C_x_PM_NOR3_X2__A3_c3 VSS N_A3_M3_g 5.91756e-17
R_x_PM_NOR3_X2__A3_r4 x_PM_NOR3_X2__A3_18 x_PM_NOR3_X2__A3_11 4.74714
R_x_PM_NOR3_X2__A3_r5 x_PM_NOR3_X2__A3_17 x_PM_NOR3_X2__A3_11 4.74714
R_x_PM_NOR3_X2__A3_r6 x_PM_NOR3_X2__A3_11 x_PM_NOR3_X2__A3_9 25.0012
R_x_PM_NOR3_X2__A3_r7 A3 x_PM_NOR3_X2__A3_9 0.2204
R_x_PM_NOR3_X2__A3_r8 N_A3_M0_g x_PM_NOR3_X2__A3_18 49.14
R_x_PM_NOR3_X2__A3_r9 N_A3_M3_g x_PM_NOR3_X2__A3_17 74.88
C_x_PM_NOR3_X2__Zalp1_c0 VSS x_PM_NOR3_X2__Zalp1_22 2.56413e-18
C_x_PM_NOR3_X2__Zalp1_c1 VSS Zalp1 5.06951e-17
C_x_PM_NOR3_X2__Zalp1_c2 VSS N_Zalp1_M2_d 2.75881e-17
C_x_PM_NOR3_X2__Zalp1_c3 VSS x_PM_NOR3_X2__Zalp1_14 6.25994e-18
C_x_PM_NOR3_X2__Zalp1_c4 VSS N_Zalp1_M5_d 2.52851e-17
C_x_PM_NOR3_X2__Zalp1_c5 VSS x_PM_NOR3_X2__Zalp1_9 8.16416e-18
C_x_PM_NOR3_X2__Zalp1_c6 VSS x_PM_NOR3_X2__Zalp1_8 4.12951e-17
C_x_PM_NOR3_X2__Zalp1_c7 VSS N_Zalp1_M3_d 2.15312e-17
R_x_PM_NOR3_X2__Zalp1_r8 Zalp1 x_PM_NOR3_X2__Zalp1_19 1.46571
R_x_PM_NOR3_X2__Zalp1_r9 x_PM_NOR3_X2__Zalp1_22 x_PM_NOR3_X2__Zalp1_18 0.143785
R_x_PM_NOR3_X2__Zalp1_r10 Zalp1 x_PM_NOR3_X2__Zalp1_18 0.868571
R_x_PM_NOR3_X2__Zalp1_r11 x_PM_NOR3_X2__Zalp1_19 x_PM_NOR3_X2__Zalp1_14 0.20978
R_x_PM_NOR3_X2__Zalp1_r12 N_Zalp1_M2_d x_PM_NOR3_X2__Zalp1_14 0.686111
R_x_PM_NOR3_X2__Zalp1_r13 x_PM_NOR3_X2__Zalp1_22 x_PM_NOR3_X2__Zalp1_10 0.143785
R_x_PM_NOR3_X2__Zalp1_r14 N_Zalp1_M5_d x_PM_NOR3_X2__Zalp1_10 0.116111
R_x_PM_NOR3_X2__Zalp1_r15 x_PM_NOR3_X2__Zalp1_22 x_PM_NOR3_X2__Zalp1_8 0.0569232
R_x_PM_NOR3_X2__Zalp1_r16 x_PM_NOR3_X2__Zalp1_9 x_PM_NOR3_X2__Zalp1_8 1.65571
R_x_PM_NOR3_X2__Zalp1_r17 x_PM_NOR3_X2__Zalp1_9 x_PM_NOR3_X2__Zalp1_4 0.212317
R_x_PM_NOR3_X2__Zalp1_r18 N_Zalp1_M3_d x_PM_NOR3_X2__Zalp1_4 0.149286
C_x_PM_NOR3_X2__A2_c0 VSS x_PM_NOR3_X2__A2_11 8.98632e-18
C_x_PM_NOR3_X2__A2_c1 VSS x_PM_NOR3_X2__A2_9 8.53584e-17
C_x_PM_NOR3_X2__A2_c2 VSS N_A2_M1_g 6.12109e-17
C_x_PM_NOR3_X2__A2_c3 VSS N_A2_M4_g 6.60015e-17
R_x_PM_NOR3_X2__A2_r4 x_PM_NOR3_X2__A2_18 x_PM_NOR3_X2__A2_11 4.74714
R_x_PM_NOR3_X2__A2_r5 x_PM_NOR3_X2__A2_17 x_PM_NOR3_X2__A2_11 4.74714
R_x_PM_NOR3_X2__A2_r6 x_PM_NOR3_X2__A2_11 x_PM_NOR3_X2__A2_9 25.0012
R_x_PM_NOR3_X2__A2_r7 A2 x_PM_NOR3_X2__A2_9 0.2204
R_x_PM_NOR3_X2__A2_r8 N_A2_M1_g x_PM_NOR3_X2__A2_18 49.14
R_x_PM_NOR3_X2__A2_r9 N_A2_M4_g x_PM_NOR3_X2__A2_17 74.88
C_x_PM_NOR3_X2__A1_c0 VSS x_PM_NOR3_X2__A1_20 1.07269e-17
C_x_PM_NOR3_X2__A1_c1 VSS x_PM_NOR3_X2__A1_14 4.59258e-17
C_x_PM_NOR3_X2__A1_c2 VSS x_PM_NOR3_X2__A1_9 3.45973e-17
C_x_PM_NOR3_X2__A1_c3 VSS N_A1_M2_g 7.00434e-17
C_x_PM_NOR3_X2__A1_c4 VSS N_A1_M5_g 6.63408e-17
R_x_PM_NOR3_X2__A1_r5 x_PM_NOR3_X2__A1_20 x_PM_NOR3_X2__A1_16 2.34
R_x_PM_NOR3_X2__A1_r6 x_PM_NOR3_X2__A1_16 x_PM_NOR3_X2__A1_14 25.0012
R_x_PM_NOR3_X2__A1_r7 x_PM_NOR3_X2__A1_14 x_PM_NOR3_X2__A1_12 0.147778
R_x_PM_NOR3_X2__A1_r8 x_PM_NOR3_X2__A1_12 x_PM_NOR3_X2__A1_9 0.095
R_x_PM_NOR3_X2__A1_r9 A1 x_PM_NOR3_X2__A1_9 0.298571
R_x_PM_NOR3_X2__A1_r10 x_PM_NOR3_X2__A1_20 x_PM_NOR3_X2__A1_5 1.95
R_x_PM_NOR3_X2__A1_r11 N_A1_M2_g x_PM_NOR3_X2__A1_5 56.94
R_x_PM_NOR3_X2__A1_r12 x_PM_NOR3_X2__A1_20 x_PM_NOR3_X2__A1_VSS 1.95
R_x_PM_NOR3_X2__A1_r13 N_A1_M5_g x_PM_NOR3_X2__A1_VSS 67.08

********************************************NOR2_X2****************************************************
M2_M2 62 N2_A5_M0_g N2_VDD_M0_s VDD PMOS_VTL W=0.390000U AS=0.040950P AD=0.054600P PS=0.990000U PD=1.060000U
M2_M3 N2_Zalp2_M1_d N2_A4_M1_g 62 VDD PMOS_VTL W=0.390000U AS=0.054600P AD=0.040950P PS=1.060000U PD=0.990000U
M2_M0 N2_Zalp2_M2_d N2_A5_M2_g N2_VSS_M2_s VSS NMOS_VTL W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M2_M1 N2_VSS_M3_d N2_A4_M3_g N2_Zalp2_M2_d VSS NMOS_VTL W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_NOR2_X2__VSS_c0 VSS N2_VSS_M3_d 1.9003e-17
C_x_PM_NOR2_X2__VSS_c1 VSS x_PM_NOR2_X2__VSS_8 1.14613e-17
C_x_PM_NOR2_X2__VSS_c2 VSS x_PM_NOR2_X2__VSS_7 5.12113e-17
C_x_PM_NOR2_X2__VSS_c3 VSS N2_VSS_M2_s 1.7976e-17
R_x_PM_NOR2_X2__VSS_r4 N2_VSS_M3_d x_PM_NOR2_X2__VSS_11 0.230714
R_x_PM_NOR2_X2__VSS_r5 VSS x_PM_NOR2_X2__VSS_8 0.357647
R_x_PM_NOR2_X2__VSS_r6 x_PM_NOR2_X2__VSS_11 x_PM_NOR2_X2__VSS_7 0.264221
R_x_PM_NOR2_X2__VSS_r7 VSS x_PM_NOR2_X2__VSS_7 0.324118
R_x_PM_NOR2_X2__VSS_r8 x_PM_NOR2_X2__VSS_8 x_PM_NOR2_X2__VSS_3 0.264221
R_x_PM_NOR2_X2__VSS_r9 N2_VSS_M2_s x_PM_NOR2_X2__VSS_3 0.230714
C_x_PM_NOR2_X2__VDD_c0 VSS VDD 5.55967e-17
C_x_PM_NOR2_X2__VDD_c1 VSS N2_VDD_M0_s 2.30938e-17
R_x_PM_NOR2_X2__VDD_r2 x_PM_NOR2_X2__VDD_10 VDD 0.0881799
R_x_PM_NOR2_X2__VDD_r3 N2_VDD_M0_s x_PM_NOR2_X2__VDD_10 0.230714
C_x_PM_NOR2_X2__A5_c0 VSS x_PM_NOR2_X2__A5_18 8.24826e-18
C_x_PM_NOR2_X2__A5_c1 VSS x_PM_NOR2_X2__A5_12 4.45792e-17
C_x_PM_NOR2_X2__A5_c2 VSS N2_A5_M0_g 9.21574e-17
C_x_PM_NOR2_X2__A5_c3 VSS N2_A5_M2_g 3.09335e-17
R_x_PM_NOR2_X2__A5_r4 x_PM_NOR2_X2__A5_18 x_PM_NOR2_X2__A5_14 3.38
R_x_PM_NOR2_X2__A5_r5 x_PM_NOR2_X2__A5_14 x_PM_NOR2_X2__A5_12 25.0012
R_x_PM_NOR2_X2__A5_r6 x_PM_NOR2_X2__A5_12 A5 0.15069
R_x_PM_NOR2_X2__A5_r7 x_PM_NOR2_X2__A5_18 x_PM_NOR2_X2__A5_5 1.95
R_x_PM_NOR2_X2__A5_r8 N2_A5_M0_g x_PM_NOR2_X2__A5_5 112.32
R_x_PM_NOR2_X2__A5_r9 x_PM_NOR2_X2__A5_18 x_PM_NOR2_X2__A5_VSS 1.95
R_x_PM_NOR2_X2__A5_r10 N2_A5_M2_g x_PM_NOR2_X2__A5_VSS 21.84
C_x_PM_NOR2_X2__Zalp2_c0 VSS N2_Zalp2_M1_d 5.96075e-17
C_x_PM_NOR2_X2__Zalp2_c1 VSS x_PM_NOR2_X2__Zalp2_9 3.74417e-17
C_x_PM_NOR2_X2__Zalp2_c2 VSS Zalp2 7.19517e-18
C_x_PM_NOR2_X2__Zalp2_c3 VSS N2_Zalp2_M2_d 8.47483e-17
R_x_PM_NOR2_X2__Zalp2_r4 N2_Zalp2_M1_d x_PM_NOR2_X2__Zalp2_11 2.91786
R_x_PM_NOR2_X2__Zalp2_r5 x_PM_NOR2_X2__Zalp2_11 x_PM_NOR2_X2__Zalp2_9 0.212317
R_x_PM_NOR2_X2__Zalp2_r6 x_PM_NOR2_X2__Zalp2_10 x_PM_NOR2_X2__Zalp2_9 0.597143
R_x_PM_NOR2_X2__Zalp2_r7 x_PM_NOR2_X2__Zalp2_10 Zalp2 0.212317
R_x_PM_NOR2_X2__Zalp2_r8 Zalp2 x_PM_NOR2_X2__Zalp2_7 0.000542857
R_x_PM_NOR2_X2__Zalp2_r9 x_PM_NOR2_X2__Zalp2_7 N2_Zalp2_M2_d 1.39731
C_x_PM_NOR2_X2__A4_c0 VSS A4 6.50458e-17
C_x_PM_NOR2_X2__A4_c1 VSS x_PM_NOR2_X2__A4_11 9.81933e-18
C_x_PM_NOR2_X2__A4_c2 VSS N2_A4_M1_g 1.07185e-16
C_x_PM_NOR2_X2__A4_c3 VSS N2_A4_M3_g 3.09279e-17
R_x_PM_NOR2_X2__A4_r4 x_PM_NOR2_X2__A4_11 x_PM_NOR2_X2__A4_16 4.42
R_x_PM_NOR2_X2__A4_r5 x_PM_NOR2_X2__A4_11 x_PM_NOR2_X2__A4_9 25.0012
R_x_PM_NOR2_X2__A4_r6 A4 x_PM_NOR2_X2__A4_9 0.15069
R_x_PM_NOR2_X2__A4_r7 x_PM_NOR2_X2__A4_16 x_PM_NOR2_X2__A4_5 1.95
R_x_PM_NOR2_X2__A4_r8 N2_A4_M1_g x_PM_NOR2_X2__A4_5 112.32
R_x_PM_NOR2_X2__A4_r9 x_PM_NOR2_X2__A4_16 x_PM_NOR2_X2__A4_VSS 1.95
R_x_PM_NOR2_X2__A4_r10 N2_A4_M3_g x_PM_NOR2_X2__A4_VSS 21.84

********************************************NAND2_X2**************************************************
M3_M2 N3_ZN3_M0_d N3_Zalp2_M0_g N3_VDD_M0_s VDD PMOS_VTL W=0.270000U AS=0.028350P AD=0.037800P PS=0.750000U PD=0.820000U
M3_M3 N3_VDD_M1_d N3_Zalp1_M1_g N3_ZN3_M0_d VDD PMOS_VTL W=0.270000U AS=0.037800P AD=0.028350P PS=0.820000U PD=0.750000U
M3_M0 63 N3_Zalp2_M2_g N3_VSS_M2_s VSS NMOS_VTL W=0.260000U AS=0.027300P AD=0.036400P PS=0.730000U PD=0.800000U
M3_M1 N3_ZN3_M3_d N3_Zalp1_M3_g 63 VSS NMOS_VTL W=0.260000U AS=0.036400P AD=0.027300P PS=0.800000U PD=0.730000U
C_x_PM_NAND2_X2__VSS_c0 VSS VSS 5.03826e-17
C_x_PM_NAND2_X2__VSS_c1 VSS x_PM_NAND2_X2__VSS_6 1.04465e-17
C_x_PM_NAND2_X2__VSS_c2 VSS N3_VSS_M2_s 1.83058e-17
R_x_PM_NAND2_X2__VSS_r3 VSS x_PM_NAND2_X2__VSS_6 0.391176
R_x_PM_NAND2_X2__VSS_r4 x_PM_NAND2_X2__VSS_6 x_PM_NAND2_X2__VSS_2 0.264221
R_x_PM_NAND2_X2__VSS_r5 N3_VSS_M2_s x_PM_NAND2_X2__VSS_2 0.230714
C_x_PM_NAND2_X2__VDD_c0 VSS N3_VDD_M1_d 4.75732e-17
C_x_PM_NAND2_X2__VDD_c1 VSS x_PM_NAND2_X2__VDD_7 4.67275e-17
C_x_PM_NAND2_X2__VDD_c2 VSS N3_VDD_M0_s 2.99432e-17
C_x_PM_NAND2_X2__VDD_c3 VSS x_PM_NAND2_X2__VDD_3 1.06496e-17
R_x_PM_NAND2_X2__VDD_r4 N3_VDD_M1_d x_PM_NAND2_X2__VDD_9 0.420714
R_x_PM_NAND2_X2__VDD_r5 VDD x_PM_NAND2_X2__VDD_8 0.195294
R_x_PM_NAND2_X2__VDD_r6 x_PM_NAND2_X2__VDD_9 x_PM_NAND2_X2__VDD_7 0.264221
R_x_PM_NAND2_X2__VDD_r7 x_PM_NAND2_X2__VDD_8 x_PM_NAND2_X2__VDD_7 0.681765
R_x_PM_NAND2_X2__VDD_r8 VDD x_PM_NAND2_X2__VDD_3 0.0689273
R_x_PM_NAND2_X2__VDD_r9 N3_VDD_M0_s x_PM_NAND2_X2__VDD_3 0.420714
C_x_PM_NAND2_X2__Zalp2_c0 VSS x_PM_NAND2_X2__Zalp2_14 7.51478e-18
C_x_PM_NAND2_X2__Zalp2_c1 VSS Zalp2 6.01437e-17
C_x_PM_NAND2_X2__Zalp2_c2 VSS N3_Zalp2_M0_g 8.26414e-17
C_x_PM_NAND2_X2__Zalp2_c3 VSS N3_Zalp2_M2_g 3.58741e-17
R_x_PM_NAND2_X2__Zalp2_r4 x_PM_NAND2_X2__Zalp2_18 x_PM_NAND2_X2__Zalp2_14 4.74714
R_x_PM_NAND2_X2__Zalp2_r5 x_PM_NAND2_X2__Zalp2_17 x_PM_NAND2_X2__Zalp2_14 4.74714
R_x_PM_NAND2_X2__Zalp2_r6 x_PM_NAND2_X2__Zalp2_14 x_PM_NAND2_X2__Zalp2_12 25.0012
R_x_PM_NAND2_X2__Zalp2_r7 x_PM_NAND2_X2__Zalp2_12 Zalp2 0.266
R_x_PM_NAND2_X2__Zalp2_r8 N3_Zalp2_M0_g x_PM_NAND2_X2__Zalp2_18 103.74
R_x_PM_NAND2_X2__Zalp2_r9 N3_Zalp2_M2_g x_PM_NAND2_X2__Zalp2_17 28.08
C_x_PM_NAND2_X2__ZN3_c0 VSS N3_ZN3_M3_d 9.46701e-17
C_x_PM_NAND2_X2__ZN3_c1 VSS x_PM_NAND2_X2__ZN3_8 7.68686e-18
C_x_PM_NAND2_X2__ZN3_c2 VSS x_PM_NAND2_X2__ZN3_7 3.24105e-17
C_x_PM_NAND2_X2__ZN3_c3 VSS N3_ZN3_M0_d 6.2878e-17
R_x_PM_NAND2_X2__ZN3_r4 ZN N3_ZN3_M3_d 1.93167
R_x_PM_NAND2_X2__ZN3_r5 ZN x_PM_NAND2_X2__ZN3_9 0.527778
R_x_PM_NAND2_X2__ZN3_r6 x_PM_NAND2_X2__ZN3_9 x_PM_NAND2_X2__ZN3_7 0.21666
R_x_PM_NAND2_X2__ZN3_r7 x_PM_NAND2_X2__ZN3_8 x_PM_NAND2_X2__ZN3_7 0.624286
R_x_PM_NAND2_X2__ZN3_r8 x_PM_NAND2_X2__ZN3_8 x_PM_NAND2_X2__ZN3_3 0.212317
R_x_PM_NAND2_X2__ZN3_r9 N3_ZN3_M0_d x_PM_NAND2_X2__ZN3_3 1.18071
C_x_PM_NAND2_X2__Zalp1_c0 VSS x_PM_NAND2_X2__Zalp1_18 1.23667e-17
C_x_PM_NAND2_X2__Zalp1_c1 VSS Zalp1 8.87208e-17
C_x_PM_NAND2_X2__Zalp1_c2 VSS N3_Zalp1_M1_g 9.96411e-17
C_x_PM_NAND2_X2__Zalp1_c3 VSS N3_Zalp1_M3_g 3.7962e-17
R_x_PM_NAND2_X2__Zalp1_r4 x_PM_NAND2_X2__Zalp1_18 x_PM_NAND2_X2__Zalp1_14 3.9
R_x_PM_NAND2_X2__Zalp1_r5 x_PM_NAND2_X2__Zalp1_14 x_PM_NAND2_X2__Zalp1_12 25.0012
R_x_PM_NAND2_X2__Zalp1_r6 x_PM_NAND2_X2__Zalp1_12 Zalp1 0.316667
R_x_PM_NAND2_X2__Zalp1_r7 x_PM_NAND2_X2__Zalp1_18 x_PM_NAND2_X2__Zalp1_5 1.95
R_x_PM_NAND2_X2__Zalp1_r8 N3_Zalp1_M1_g x_PM_NAND2_X2__Zalp1_5 103.74
R_x_PM_NAND2_X2__Zalp1_r9 x_PM_NAND2_X2__Zalp1_18 x_PM_NAND2_X2__Zalp1_VSS 1.95
R_x_PM_NAND2_X2__Zalp1_r10 N3_Zalp1_M3_g x_PM_NAND2_X2__Zalp1_VSS 28.08
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
