.SUBCKT or3 A1 A2 A3 VDD VSS ZN 
M_M4 8 N_A1_M0_g N_3_M0_s VDD PMOS_VTL L=0.050U W=0.260000U AS=0.027300P AD=0.036400P PS=0.730000U PD=0.800000U
M_M5 9 N_A2_M1_g 8 VDD PMOS_VTL L=0.050U W=0.260000U AS=0.036400P AD=0.036400P PS=0.800000U PD=0.800000U
M_M6 N_VDD_M2_d N_A3_M2_g 9 VDD PMOS_VTL L=0.050U W=0.260000U AS=0.036400P AD=0.037300P PS=0.800000U PD=0.820000U
M_M7 N_ZN_M3_d N_3_M3_g N_VDD_M2_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037300P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 N_VSS_M4_d N_A1_M4_g N_3_M4_s VSS NMOS_VTL L=0.050U W=0.090000U AS=0.009450P AD=0.012600P PS=0.390000U PD=0.460000U
M_M1 N_3_M5_d N_A2_M5_g N_VSS_M4_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.012600P PS=0.460000U PD=0.460000U
M_M2 N_VSS_M6_d N_A3_M6_g N_3_M5_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.020700P PS=0.460000U PD=0.640000U
M_M3 N_ZN_M7_d N_3_M7_g N_VSS_M6_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.020700P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_OR3_X2__VSS_c0 VSS x_PM_OR3_X2__VSS_20 3.00757e-17
C_x_PM_OR3_X2__VSS_c1 VSS x_PM_OR3_X2__VSS_19 4.32297e-17
C_x_PM_OR3_X2__VSS_c2 VSS N_VSS_M6_d 3.4177e-17
C_x_PM_OR3_X2__VSS_c3 VSS x_PM_OR3_X2__VSS_9 3.33766e-17
C_x_PM_OR3_X2__VSS_c4 VSS N_VSS_M4_d 3.48682e-17
R_x_PM_OR3_X2__VSS_r5 x_PM_OR3_X2__VSS_20 x_PM_OR3_X2__VSS_13 0.145286
R_x_PM_OR3_X2__VSS_r6 N_VSS_M6_d x_PM_OR3_X2__VSS_13 0.637857
R_x_PM_OR3_X2__VSS_r7 x_PM_OR3_X2__VSS_19 x_PM_OR3_X2__VSS_10 0.0731438
R_x_PM_OR3_X2__VSS_r8 VSS x_PM_OR3_X2__VSS_10 0.346471
R_x_PM_OR3_X2__VSS_r9 x_PM_OR3_X2__VSS_20 x_PM_OR3_X2__VSS_9 0.0731438
R_x_PM_OR3_X2__VSS_r10 VSS x_PM_OR3_X2__VSS_9 0.346471
R_x_PM_OR3_X2__VSS_r11 x_PM_OR3_X2__VSS_19 x_PM_OR3_X2__VSS_5 0.145286
R_x_PM_OR3_X2__VSS_r12 N_VSS_M4_d x_PM_OR3_X2__VSS_5 0.637857
C_x_PM_OR3_X2__VDD_c0 VSS x_PM_OR3_X2__VDD_12 2.99573e-17
C_x_PM_OR3_X2__VDD_c1 VSS N_VDD_M2_d 2.4519e-17
C_x_PM_OR3_X2__VDD_c2 VSS x_PM_OR3_X2__VDD_2 6.11137e-17
R_x_PM_OR3_X2__VDD_r3 x_PM_OR3_X2__VDD_12 x_PM_OR3_X2__VDD_6 0.145286
R_x_PM_OR3_X2__VDD_r4 N_VDD_M2_d x_PM_OR3_X2__VDD_6 0.230714
R_x_PM_OR3_X2__VDD_r5 x_PM_OR3_X2__VDD_12 x_PM_OR3_X2__VDD_2 0.0731438
R_x_PM_OR3_X2__VDD_r6 VDD x_PM_OR3_X2__VDD_2 0.346471
C_x_PM_OR3_X2__3_c0 VSS x_PM_OR3_X2__3_36 1.25891e-17
C_x_PM_OR3_X2__3_c1 VSS x_PM_OR3_X2__3_28 3.72813e-17
C_x_PM_OR3_X2__3_c2 VSS x_PM_OR3_X2__3_27 6.83849e-18
C_x_PM_OR3_X2__3_c3 VSS N_3_M0_s 1.93365e-17
C_x_PM_OR3_X2__3_c4 VSS x_PM_OR3_X2__3_22 2.78594e-18
C_x_PM_OR3_X2__3_c5 VSS x_PM_OR3_X2__3_20 1.68546e-17
C_x_PM_OR3_X2__3_c6 VSS x_PM_OR3_X2__3_19 4.72915e-17
C_x_PM_OR3_X2__3_c7 VSS x_PM_OR3_X2__3_16 4.23999e-17
C_x_PM_OR3_X2__3_c8 VSS x_PM_OR3_X2__3_15 5.85797e-17
C_x_PM_OR3_X2__3_c9 VSS x_PM_OR3_X2__3_13 4.65821e-17
C_x_PM_OR3_X2__3_c10 VSS N_3_M3_g 9.93078e-17
C_x_PM_OR3_X2__3_c11 VSS N_3_M7_g 3.18899e-17
R_x_PM_OR3_X2__3_r12 x_PM_OR3_X2__3_36 x_PM_OR3_X2__3_34 4.42
R_x_PM_OR3_X2__3_r13 x_PM_OR3_X2__3_34 x_PM_OR3_X2__3_31 25.0012
R_x_PM_OR3_X2__3_r14 x_PM_OR3_X2__3_31 x_PM_OR3_X2__3_28 0.176429
R_x_PM_OR3_X2__3_r15 x_PM_OR3_X2__3_27 x_PM_OR3_X2__3_21 0.179556
R_x_PM_OR3_X2__3_r16 x_PM_OR3_X2__3_28 x_PM_OR3_X2__3_20 0.095
R_x_PM_OR3_X2__3_r17 x_PM_OR3_X2__3_21 x_PM_OR3_X2__3_20 0.868571
R_x_PM_OR3_X2__3_r18 x_PM_OR3_X2__3_27 x_PM_OR3_X2__3_19 0.026987
R_x_PM_OR3_X2__3_r19 x_PM_OR3_X2__3_19 N_3_M5_d 0.548724
R_x_PM_OR3_X2__3_r20 x_PM_OR3_X2__3_22 x_PM_OR3_X2__3_17 0.0604376
R_x_PM_OR3_X2__3_r21 x_PM_OR3_X2__3_27 x_PM_OR3_X2__3_16 0.179556
R_x_PM_OR3_X2__3_r22 x_PM_OR3_X2__3_17 x_PM_OR3_X2__3_16 1.68286
R_x_PM_OR3_X2__3_r23 x_PM_OR3_X2__3_15 N_3_M0_s 0.297071
R_x_PM_OR3_X2__3_r24 x_PM_OR3_X2__3_22 x_PM_OR3_X2__3_14 0.140052
R_x_PM_OR3_X2__3_r25 x_PM_OR3_X2__3_15 x_PM_OR3_X2__3_14 3.17571
R_x_PM_OR3_X2__3_r26 x_PM_OR3_X2__3_22 x_PM_OR3_X2__3_13 0.140052
R_x_PM_OR3_X2__3_r27 x_PM_OR3_X2__3_13 N_3_M4_s 0.467567
R_x_PM_OR3_X2__3_r28 x_PM_OR3_X2__3_36 x_PM_OR3_X2__3_5 1.95
R_x_PM_OR3_X2__3_r29 N_3_M3_g x_PM_OR3_X2__3_5 109.98
R_x_PM_OR3_X2__3_r30 x_PM_OR3_X2__3_36 x_PM_OR3_X2__3_VSS 1.95
R_x_PM_OR3_X2__3_r31 N_3_M7_g x_PM_OR3_X2__3_VSS 21.84
C_x_PM_OR3_X2__A1_c0 VSS A1 6.85526e-17
C_x_PM_OR3_X2__A1_c1 VSS x_PM_OR3_X2__A1_11 9.92086e-18
C_x_PM_OR3_X2__A1_c2 VSS N_A1_M0_g 7.53703e-17
C_x_PM_OR3_X2__A1_c3 VSS N_A1_M4_g 5.78093e-17
R_x_PM_OR3_X2__A1_r4 x_PM_OR3_X2__A1_18 x_PM_OR3_X2__A1_11 4.7687
R_x_PM_OR3_X2__A1_r5 x_PM_OR3_X2__A1_17 x_PM_OR3_X2__A1_11 4.7687
R_x_PM_OR3_X2__A1_r6 x_PM_OR3_X2__A1_11 x_PM_OR3_X2__A1_9 25.0012
R_x_PM_OR3_X2__A1_r7 A1 x_PM_OR3_X2__A1_9 0.210357
R_x_PM_OR3_X2__A1_r8 N_A1_M0_g x_PM_OR3_X2__A1_18 80.34
R_x_PM_OR3_X2__A1_r9 N_A1_M4_g x_PM_OR3_X2__A1_17 59.28
C_x_PM_OR3_X2__A2_c0 VSS A2 4.50716e-17
C_x_PM_OR3_X2__A2_c1 VSS x_PM_OR3_X2__A2_11 1.07434e-17
C_x_PM_OR3_X2__A2_c2 VSS N_A2_M1_g 6.86698e-17
C_x_PM_OR3_X2__A2_c3 VSS N_A2_M5_g 5.1379e-17
R_x_PM_OR3_X2__A2_r4 x_PM_OR3_X2__A2_11 x_PM_OR3_X2__A2_16 3.38
R_x_PM_OR3_X2__A2_r5 x_PM_OR3_X2__A2_11 x_PM_OR3_X2__A2_9 25.0012
R_x_PM_OR3_X2__A2_r6 A2 x_PM_OR3_X2__A2_9 0.156071
R_x_PM_OR3_X2__A2_r7 x_PM_OR3_X2__A2_16 x_PM_OR3_X2__A2_5 1.95
R_x_PM_OR3_X2__A2_r8 N_A2_M1_g x_PM_OR3_X2__A2_5 80.34
R_x_PM_OR3_X2__A2_r9 x_PM_OR3_X2__A2_16 x_PM_OR3_X2__A2_VSS 1.95
R_x_PM_OR3_X2__A2_r10 N_A2_M5_g x_PM_OR3_X2__A2_VSS 59.28
C_x_PM_OR3_X2__A3_c0 VSS x_PM_OR3_X2__A3_11 8.5453e-18
C_x_PM_OR3_X2__A3_c1 VSS x_PM_OR3_X2__A3_9 4.53477e-17
C_x_PM_OR3_X2__A3_c2 VSS N_A3_M2_g 3.69294e-17
C_x_PM_OR3_X2__A3_c3 VSS N_A3_M6_g 8.38994e-17
R_x_PM_OR3_X2__A3_r4 x_PM_OR3_X2__A3_16 x_PM_OR3_X2__A3_11 4.7687
R_x_PM_OR3_X2__A3_r5 x_PM_OR3_X2__A3_15 x_PM_OR3_X2__A3_11 4.7687
R_x_PM_OR3_X2__A3_r6 x_PM_OR3_X2__A3_11 x_PM_OR3_X2__A3_9 25.0012
R_x_PM_OR3_X2__A3_r7 A3 x_PM_OR3_X2__A3_9 0.226453
R_x_PM_OR3_X2__A3_r8 N_A3_M2_g x_PM_OR3_X2__A3_16 28.08
R_x_PM_OR3_X2__A3_r9 N_A3_M6_g x_PM_OR3_X2__A3_15 111.54
C_x_PM_OR3_X2__ZN_c0 VSS N_ZN_M7_d 1.0669e-16
R_x_PM_OR3_X2__ZN_r1 N_ZN_M3_d ZN 2.42929
R_x_PM_OR3_X2__ZN_r2 ZN N_ZN_M7_d 1.75071
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
