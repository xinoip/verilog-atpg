.SUBCKT and4 A1 A2 A3 A4 VDD VSS ZN 
M_M5 N_3_M0_d N_A1_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.135000U  AS=0.014175P AD=0.018900P PS=0.480000U PD=0.550000U
M_M6 N_VDD_M1_d N_A2_M1_g N_3_M0_d VDD PMOS_VTL L=0.050U W=0.135000U  AS=0.018900P AD=0.018900P PS=0.550000U PD=0.550000U
M_M7 N_3_M2_d N_A3_M2_g N_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.135000U  AS=0.018900P AD=0.018900P PS=0.550000U PD=0.550000U
M_M8 N_VDD_M3_d N_A4_M3_g N_3_M2_d VDD PMOS_VTL L=0.050U W=0.135000U  AS=0.018900P AD=0.028350P PS=0.550000U PD=0.820000U
M_M9 N_ZN_M4_d N_3_M4_g N_VDD_M3_d VDD PMOS_VTL L=0.050U W=0.270000U  AS=0.028350P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 9 N_A1_M5_g N_3_M5_s VSS NMOS_VTL L=0.050U W=0.215000U  AS=0.022575P AD=0.030100P PS=0.640000U PD=0.710000U
M_M1 10 N_A2_M6_g 9 VSS NMOS_VTL L=0.050U W=0.215000U  AS=0.030100P AD=0.030100P PS=0.710000U PD=0.710000U
M_M2 11 N_A3_M7_g 10 VSS NMOS_VTL L=0.050U W=0.215000U  AS=0.030100P AD=0.030100P PS=0.710000U PD=0.710000U
M_M3 N_VSS_M8_d N_A4_M8_g 11 VSS NMOS_VTL L=0.050U W=0.215000U  AS=0.030100P AD=0.027650P PS=0.710000U PD=0.710000U
M_M4 N_ZN_M9_d N_3_M9_g N_VSS_M8_d VSS NMOS_VTL L=0.050U W=0.180000U  AS=0.027650P AD=0.018900P PS=0.710000U PD=0.570000U
C_x_PM_AND4_X2__VSS_c0 VSS x_PM_AND4_X2__VSS_12 4.48532e-17
C_x_PM_AND4_X2__VSS_c1 VSS N_VSS_M8_d 2.45741e-17
C_x_PM_AND4_X2__VSS_c2 VSS x_PM_AND4_X2__VSS_2 9.14419e-17
R_x_PM_AND4_X2__VSS_r3 x_PM_AND4_X2__VSS_12 x_PM_AND4_X2__VSS_6 0.145286
R_x_PM_AND4_X2__VSS_r4 N_VSS_M8_d x_PM_AND4_X2__VSS_6 0.230714
R_x_PM_AND4_X2__VSS_r5 x_PM_AND4_X2__VSS_12 x_PM_AND4_X2__VSS_2 0.0731438
R_x_PM_AND4_X2__VSS_r6 VSS x_PM_AND4_X2__VSS_2 0.502941
C_x_PM_AND4_X2__VDD_c0 VSS x_PM_AND4_X2__VDD_25 4.45927e-17
C_x_PM_AND4_X2__VDD_c1 VSS x_PM_AND4_X2__VDD_24 2.84978e-18
C_x_PM_AND4_X2__VDD_c2 VSS N_VDD_M3_d 2.75841e-17
C_x_PM_AND4_X2__VDD_c3 VSS x_PM_AND4_X2__VDD_14 3.21954e-17
C_x_PM_AND4_X2__VDD_c4 VSS N_VDD_M1_d 2.5303e-17
C_x_PM_AND4_X2__VDD_c5 VSS x_PM_AND4_X2__VDD_9 1.08478e-17
C_x_PM_AND4_X2__VDD_c6 VSS x_PM_AND4_X2__VDD_8 3.13029e-17
C_x_PM_AND4_X2__VDD_c7 VSS N_VDD_M0_s 1.41211e-17
R_x_PM_AND4_X2__VDD_r8 x_PM_AND4_X2__VDD_25 x_PM_AND4_X2__VDD_18 0.145286
R_x_PM_AND4_X2__VDD_r9 N_VDD_M3_d x_PM_AND4_X2__VDD_18 0.420714
R_x_PM_AND4_X2__VDD_r10 x_PM_AND4_X2__VDD_24 x_PM_AND4_X2__VDD_15 0.0731438
R_x_PM_AND4_X2__VDD_r11 VDD x_PM_AND4_X2__VDD_15 0.19
R_x_PM_AND4_X2__VDD_r12 x_PM_AND4_X2__VDD_25 x_PM_AND4_X2__VDD_14 0.0731438
R_x_PM_AND4_X2__VDD_r13 VDD x_PM_AND4_X2__VDD_14 0.502941
R_x_PM_AND4_X2__VDD_r14 x_PM_AND4_X2__VDD_24 x_PM_AND4_X2__VDD_10 0.145286
R_x_PM_AND4_X2__VDD_r15 N_VDD_M1_d x_PM_AND4_X2__VDD_10 0.420714
R_x_PM_AND4_X2__VDD_r16 x_PM_AND4_X2__VDD_24 x_PM_AND4_X2__VDD_8 0.0731438
R_x_PM_AND4_X2__VDD_r17 x_PM_AND4_X2__VDD_9 x_PM_AND4_X2__VDD_8 0.681765
R_x_PM_AND4_X2__VDD_r18 x_PM_AND4_X2__VDD_9 x_PM_AND4_X2__VDD_4 0.264221
R_x_PM_AND4_X2__VDD_r19 N_VDD_M0_s x_PM_AND4_X2__VDD_4 0.420714
C_x_PM_AND4_X2__3_c0 VSS x_PM_AND4_X2__3_40 1.12164e-17
C_x_PM_AND4_X2__3_c1 VSS x_PM_AND4_X2__3_33 2.06085e-18
C_x_PM_AND4_X2__3_c2 VSS N_3_M5_s 2.68504e-17
C_x_PM_AND4_X2__3_c3 VSS x_PM_AND4_X2__3_27 8.75385e-17
C_x_PM_AND4_X2__3_c4 VSS x_PM_AND4_X2__3_26 5.12014e-17
C_x_PM_AND4_X2__3_c5 VSS x_PM_AND4_X2__3_24 3.28897e-17
C_x_PM_AND4_X2__3_c6 VSS N_3_M2_d 3.41478e-17
C_x_PM_AND4_X2__3_c7 VSS x_PM_AND4_X2__3_19 1.0345e-17
C_x_PM_AND4_X2__3_c8 VSS x_PM_AND4_X2__3_18 2.94817e-17
C_x_PM_AND4_X2__3_c9 VSS N_3_M0_d 3.60348e-17
C_x_PM_AND4_X2__3_c10 VSS x_PM_AND4_X2__3_12 1.17003e-16
C_x_PM_AND4_X2__3_c11 VSS N_3_M4_g 1.01497e-16
C_x_PM_AND4_X2__3_c12 VSS N_3_M9_g 3.57135e-17
R_x_PM_AND4_X2__3_r13 x_PM_AND4_X2__3_40 x_PM_AND4_X2__3_38 3.38
R_x_PM_AND4_X2__3_r14 x_PM_AND4_X2__3_38 x_PM_AND4_X2__3_36 25.0012
R_x_PM_AND4_X2__3_r15 x_PM_AND4_X2__3_36 x_PM_AND4_X2__3_34 0.259615
R_x_PM_AND4_X2__3_r16 x_PM_AND4_X2__3_31 N_3_M5_s 0.285
R_x_PM_AND4_X2__3_r17 x_PM_AND4_X2__3_36 x_PM_AND4_X2__3_26 0.292415
R_x_PM_AND4_X2__3_r18 x_PM_AND4_X2__3_27 x_PM_AND4_X2__3_26 2.93143
R_x_PM_AND4_X2__3_r19 x_PM_AND4_X2__3_33 x_PM_AND4_X2__3_25 0.160909
R_x_PM_AND4_X2__3_r20 x_PM_AND4_X2__3_27 x_PM_AND4_X2__3_24 0.212317
R_x_PM_AND4_X2__3_r21 x_PM_AND4_X2__3_25 x_PM_AND4_X2__3_24 0.787143
R_x_PM_AND4_X2__3_r22 x_PM_AND4_X2__3_33 x_PM_AND4_X2__3_20 0.0418175
R_x_PM_AND4_X2__3_r23 N_3_M2_d x_PM_AND4_X2__3_20 0.610714
R_x_PM_AND4_X2__3_r24 x_PM_AND4_X2__3_33 x_PM_AND4_X2__3_18 0.160909
R_x_PM_AND4_X2__3_r25 x_PM_AND4_X2__3_19 x_PM_AND4_X2__3_18 1.65571
R_x_PM_AND4_X2__3_r26 x_PM_AND4_X2__3_19 x_PM_AND4_X2__3_14 0.212317
R_x_PM_AND4_X2__3_r27 N_3_M0_d x_PM_AND4_X2__3_14 0.610714
R_x_PM_AND4_X2__3_r28 x_PM_AND4_X2__3_31 x_PM_AND4_X2__3_13 0.095
R_x_PM_AND4_X2__3_r29 x_PM_AND4_X2__3_34 x_PM_AND4_X2__3_12 0.100962
R_x_PM_AND4_X2__3_r30 x_PM_AND4_X2__3_13 x_PM_AND4_X2__3_12 3.85429
R_x_PM_AND4_X2__3_r31 x_PM_AND4_X2__3_40 x_PM_AND4_X2__3_5 1.95
R_x_PM_AND4_X2__3_r32 N_3_M4_g x_PM_AND4_X2__3_5 111.54
R_x_PM_AND4_X2__3_r33 x_PM_AND4_X2__3_40 x_PM_AND4_X2__3_VSS 1.95
R_x_PM_AND4_X2__3_r34 N_3_M9_g x_PM_AND4_X2__3_VSS 26.52
C_x_PM_AND4_X2__A1_c0 VSS x_PM_AND4_X2__A1_14 7.4392e-18
C_x_PM_AND4_X2__A1_c1 VSS x_PM_AND4_X2__A1_12 4.24683e-17
C_x_PM_AND4_X2__A1_c2 VSS N_A1_M0_g 7.33374e-17
C_x_PM_AND4_X2__A1_c3 VSS N_A1_M5_g 4.39981e-17
R_x_PM_AND4_X2__A1_r4 x_PM_AND4_X2__A1_18 x_PM_AND4_X2__A1_14 4.7687
R_x_PM_AND4_X2__A1_r5 x_PM_AND4_X2__A1_17 x_PM_AND4_X2__A1_14 4.7687
R_x_PM_AND4_X2__A1_r6 x_PM_AND4_X2__A1_14 x_PM_AND4_X2__A1_12 25.0012
R_x_PM_AND4_X2__A1_r7 x_PM_AND4_X2__A1_12 A1 0.2375
R_x_PM_AND4_X2__A1_r8 N_A1_M0_g x_PM_AND4_X2__A1_18 106.47
R_x_PM_AND4_X2__A1_r9 N_A1_M5_g x_PM_AND4_X2__A1_17 39.39
C_x_PM_AND4_X2__A2_c0 VSS x_PM_AND4_X2__A2_14 8.42144e-18
C_x_PM_AND4_X2__A2_c1 VSS x_PM_AND4_X2__A2_12 2.222e-17
C_x_PM_AND4_X2__A2_c2 VSS N_A2_M1_g 5.45019e-17
C_x_PM_AND4_X2__A2_c3 VSS N_A2_M6_g 7.16293e-17
R_x_PM_AND4_X2__A2_r4 x_PM_AND4_X2__A2_18 x_PM_AND4_X2__A2_14 4.7687
R_x_PM_AND4_X2__A2_r5 x_PM_AND4_X2__A2_17 x_PM_AND4_X2__A2_14 4.7687
R_x_PM_AND4_X2__A2_r6 x_PM_AND4_X2__A2_14 x_PM_AND4_X2__A2_12 25.0012
R_x_PM_AND4_X2__A2_r7 x_PM_AND4_X2__A2_12 A2 0.169643
R_x_PM_AND4_X2__A2_r8 N_A2_M1_g x_PM_AND4_X2__A2_18 62.79
R_x_PM_AND4_X2__A2_r9 N_A2_M6_g x_PM_AND4_X2__A2_17 83.07
C_x_PM_AND4_X2__A3_c0 VSS x_PM_AND4_X2__A3_14 9.23042e-18
C_x_PM_AND4_X2__A3_c1 VSS x_PM_AND4_X2__A3_12 5.936e-17
C_x_PM_AND4_X2__A3_c2 VSS N_A3_M2_g 8.12259e-17
C_x_PM_AND4_X2__A3_c3 VSS N_A3_M7_g 4.54243e-17
R_x_PM_AND4_X2__A3_r4 x_PM_AND4_X2__A3_18 x_PM_AND4_X2__A3_14 4.74714
R_x_PM_AND4_X2__A3_r5 x_PM_AND4_X2__A3_17 x_PM_AND4_X2__A3_14 4.74714
R_x_PM_AND4_X2__A3_r6 x_PM_AND4_X2__A3_14 x_PM_AND4_X2__A3_12 25.0012
R_x_PM_AND4_X2__A3_r7 x_PM_AND4_X2__A3_12 A3 0.156071
R_x_PM_AND4_X2__A3_r8 N_A3_M2_g x_PM_AND4_X2__A3_18 106.47
R_x_PM_AND4_X2__A3_r9 N_A3_M7_g x_PM_AND4_X2__A3_17 39.39
C_x_PM_AND4_X2__A4_c0 VSS x_PM_AND4_X2__A4_14 8.80305e-18
C_x_PM_AND4_X2__A4_c1 VSS x_PM_AND4_X2__A4_12 8.0586e-17
C_x_PM_AND4_X2__A4_c2 VSS N_A4_M3_g 8.26834e-17
C_x_PM_AND4_X2__A4_c3 VSS N_A4_M8_g 4.63995e-17
R_x_PM_AND4_X2__A4_r4 x_PM_AND4_X2__A4_18 x_PM_AND4_X2__A4_14 4.7687
R_x_PM_AND4_X2__A4_r5 x_PM_AND4_X2__A4_17 x_PM_AND4_X2__A4_14 4.7687
R_x_PM_AND4_X2__A4_r6 x_PM_AND4_X2__A4_14 x_PM_AND4_X2__A4_12 25.0012
R_x_PM_AND4_X2__A4_r7 x_PM_AND4_X2__A4_12 A4 0.169643
R_x_PM_AND4_X2__A4_r8 N_A4_M3_g x_PM_AND4_X2__A4_18 106.47
R_x_PM_AND4_X2__A4_r9 N_A4_M8_g x_PM_AND4_X2__A4_17 39.39
C_x_PM_AND4_X2__ZN_c0 VSS N_ZN_M9_d 3.54907e-17
C_x_PM_AND4_X2__ZN_c1 VSS ZN 8.1492e-17
C_x_PM_AND4_X2__ZN_c2 VSS N_ZN_M4_d 4.91094e-17
C_x_PM_AND4_X2__ZN_c3 VSS x_PM_AND4_X2__ZN_3 6.62394e-18
R_x_PM_AND4_X2__ZN_r4 ZN x_PM_AND4_X2__ZN_8 1.87286
R_x_PM_AND4_X2__ZN_r5 x_PM_AND4_X2__ZN_7 N_ZN_M9_d 0.30478
R_x_PM_AND4_X2__ZN_r6 ZN x_PM_AND4_X2__ZN_7 1.84571
R_x_PM_AND4_X2__ZN_r7 x_PM_AND4_X2__ZN_8 x_PM_AND4_X2__ZN_3 0.20978
R_x_PM_AND4_X2__ZN_r8 N_ZN_M4_d x_PM_AND4_X2__ZN_3 0.686111
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
