.SUBCKT and3 A1 A2 A3 VDD VSS ZN 
M_M4 N_VDD_M0_d N_A1_M0_g N_3_M0_s VDD PMOS_VTL L=0.050U W=0.135000U AS=0.014175P AD=0.018900P PS=0.480000U PD=0.550000U
M_M5 N_3_M1_d N_A2_M1_g N_VDD_M0_d VDD PMOS_VTL L=0.050U W=0.135000U AS=0.018900P AD=0.018900P PS=0.550000U PD=0.550000U
M_M6 N_VDD_M2_d N_A3_M2_g N_3_M1_d VDD PMOS_VTL L=0.050U W=0.135000U AS=0.018900P AD=0.028350P PS=0.550000U PD=0.820000U
M_M7 N_ZN_M3_d N_3_M3_g N_VDD_M2_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 8 N_A1_M4_g N_3_M4_s VSS NMOS_VTL L=0.050U W=0.170000U AS=0.017850P AD=0.023800P PS=0.550000U PD=0.620000U
M_M1 9 N_A2_M5_g 8 VSS NMOS_VTL L=0.050U W=0.170000U AS=0.023800P AD=0.023800P PS=0.620000U PD=0.620000U
M_M2 N_VSS_M6_d N_A3_M6_g 9 VSS NMOS_VTL L=0.050U W=0.170000U AS=0.023800P AD=0.024700P PS=0.620000U PD=0.640000U
M_M3 N_ZN_M7_d N_3_M7_g N_VSS_M6_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.024700P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_AND3_X2__VSS_c0 VSS x_PM_AND3_X2__VSS_12 4.21405e-17
C_x_PM_AND3_X2__VSS_c1 VSS N_VSS_M6_d 2.36734e-17
C_x_PM_AND3_X2__VSS_c2 VSS x_PM_AND3_X2__VSS_2 7.71966e-17
R_x_PM_AND3_X2__VSS_r3 x_PM_AND3_X2__VSS_12 x_PM_AND3_X2__VSS_6 0.145286
R_x_PM_AND3_X2__VSS_r4 N_VSS_M6_d x_PM_AND3_X2__VSS_6 0.230714
R_x_PM_AND3_X2__VSS_r5 x_PM_AND3_X2__VSS_12 x_PM_AND3_X2__VSS_2 0.0731438
R_x_PM_AND3_X2__VSS_r6 VSS x_PM_AND3_X2__VSS_2 0.290588
C_x_PM_AND3_X2__VDD_c0 VSS x_PM_AND3_X2__VDD_20 4.53039e-17
C_x_PM_AND3_X2__VDD_c1 VSS x_PM_AND3_X2__VDD_19 3.68815e-17
C_x_PM_AND3_X2__VDD_c2 VSS N_VDD_M2_d 3.50284e-17
C_x_PM_AND3_X2__VDD_c3 VSS x_PM_AND3_X2__VDD_9 3.25732e-17
C_x_PM_AND3_X2__VDD_c4 VSS N_VDD_M0_d 3.52926e-17
R_x_PM_AND3_X2__VDD_r5 x_PM_AND3_X2__VDD_20 x_PM_AND3_X2__VDD_13 0.145286
R_x_PM_AND3_X2__VDD_r6 N_VDD_M2_d x_PM_AND3_X2__VDD_13 0.420714
R_x_PM_AND3_X2__VDD_r7 x_PM_AND3_X2__VDD_19 x_PM_AND3_X2__VDD_10 0.0731438
R_x_PM_AND3_X2__VDD_r8 VDD x_PM_AND3_X2__VDD_10 0.402353
R_x_PM_AND3_X2__VDD_r9 x_PM_AND3_X2__VDD_20 x_PM_AND3_X2__VDD_9 0.0731438
R_x_PM_AND3_X2__VDD_r10 VDD x_PM_AND3_X2__VDD_9 0.290588
R_x_PM_AND3_X2__VDD_r11 x_PM_AND3_X2__VDD_19 x_PM_AND3_X2__VDD_5 0.145286
R_x_PM_AND3_X2__VDD_r12 N_VDD_M0_d x_PM_AND3_X2__VDD_5 0.420714
C_x_PM_AND3_X2__3_c0 VSS x_PM_AND3_X2__3_44 1.14374e-17
C_x_PM_AND3_X2__3_c1 VSS x_PM_AND3_X2__3_41 1.04375e-17
C_x_PM_AND3_X2__3_c2 VSS x_PM_AND3_X2__3_40 3.30128e-17
C_x_PM_AND3_X2__3_c3 VSS x_PM_AND3_X2__3_39 3.47774e-18
C_x_PM_AND3_X2__3_c4 VSS x_PM_AND3_X2__3_38 7.12662e-17
C_x_PM_AND3_X2__3_c5 VSS x_PM_AND3_X2__3_35 9.3384e-18
C_x_PM_AND3_X2__3_c6 VSS x_PM_AND3_X2__3_32 6.87787e-18
C_x_PM_AND3_X2__3_c7 VSS x_PM_AND3_X2__3_28 4.77545e-17
C_x_PM_AND3_X2__3_c8 VSS N_3_M1_d 3.07979e-17
C_x_PM_AND3_X2__3_c9 VSS x_PM_AND3_X2__3_23 4.21984e-18
C_x_PM_AND3_X2__3_c10 VSS x_PM_AND3_X2__3_22 3.23292e-17
C_x_PM_AND3_X2__3_c11 VSS x_PM_AND3_X2__3_21 1.39555e-17
C_x_PM_AND3_X2__3_c12 VSS x_PM_AND3_X2__3_20 1.02137e-16
C_x_PM_AND3_X2__3_c13 VSS N_3_M0_s 2.59812e-17
C_x_PM_AND3_X2__3_c14 VSS N_3_M4_s 2.29228e-17
C_x_PM_AND3_X2__3_c15 VSS N_3_M3_g 7.13801e-17
C_x_PM_AND3_X2__3_c16 VSS N_3_M7_g 6.00305e-17
R_x_PM_AND3_X2__3_r17 x_PM_AND3_X2__3_44 x_PM_AND3_X2__3_42 3.38
R_x_PM_AND3_X2__3_r18 x_PM_AND3_X2__3_38 x_PM_AND3_X2__3_41 1.81857
R_x_PM_AND3_X2__3_r19 x_PM_AND3_X2__3_42 x_PM_AND3_X2__3_35 25.0012
R_x_PM_AND3_X2__3_r20 x_PM_AND3_X2__3_41 x_PM_AND3_X2__3_33 0.196927
R_x_PM_AND3_X2__3_r21 x_PM_AND3_X2__3_35 x_PM_AND3_X2__3_33 0.130625
R_x_PM_AND3_X2__3_r22 x_PM_AND3_X2__3_40 x_PM_AND3_X2__3_32 0.196927
R_x_PM_AND3_X2__3_r23 x_PM_AND3_X2__3_35 x_PM_AND3_X2__3_32 0.130625
R_x_PM_AND3_X2__3_r24 x_PM_AND3_X2__3_40 x_PM_AND3_X2__3_30 1.14
R_x_PM_AND3_X2__3_r25 x_PM_AND3_X2__3_39 x_PM_AND3_X2__3_29 0.160909
R_x_PM_AND3_X2__3_r26 x_PM_AND3_X2__3_38 x_PM_AND3_X2__3_28 0.212317
R_x_PM_AND3_X2__3_r27 x_PM_AND3_X2__3_29 x_PM_AND3_X2__3_28 0.922857
R_x_PM_AND3_X2__3_r28 x_PM_AND3_X2__3_39 x_PM_AND3_X2__3_24 0.0418175
R_x_PM_AND3_X2__3_r29 N_3_M1_d x_PM_AND3_X2__3_24 0.393571
R_x_PM_AND3_X2__3_r30 x_PM_AND3_X2__3_39 x_PM_AND3_X2__3_22 0.160909
R_x_PM_AND3_X2__3_r31 x_PM_AND3_X2__3_23 x_PM_AND3_X2__3_22 1.65571
R_x_PM_AND3_X2__3_r32 x_PM_AND3_X2__3_30 x_PM_AND3_X2__3_20 0.212317
R_x_PM_AND3_X2__3_r33 x_PM_AND3_X2__3_21 x_PM_AND3_X2__3_20 2.95857
R_x_PM_AND3_X2__3_r34 x_PM_AND3_X2__3_23 x_PM_AND3_X2__3_16 0.212317
R_x_PM_AND3_X2__3_r35 N_3_M0_s x_PM_AND3_X2__3_16 0.393571
R_x_PM_AND3_X2__3_r36 x_PM_AND3_X2__3_21 x_PM_AND3_X2__3_12 0.212317
R_x_PM_AND3_X2__3_r37 N_3_M4_s x_PM_AND3_X2__3_12 0.339286
R_x_PM_AND3_X2__3_r38 x_PM_AND3_X2__3_44 x_PM_AND3_X2__3_5 1.95
R_x_PM_AND3_X2__3_r39 N_3_M3_g x_PM_AND3_X2__3_5 73.32
R_x_PM_AND3_X2__3_r40 x_PM_AND3_X2__3_44 x_PM_AND3_X2__3_VSS 1.95
R_x_PM_AND3_X2__3_r41 N_3_M7_g x_PM_AND3_X2__3_VSS 64.74
C_x_PM_AND3_X2__A1_c0 VSS x_PM_AND3_X2__A1_14 7.47882e-18
C_x_PM_AND3_X2__A1_c1 VSS x_PM_AND3_X2__A1_12 5.57778e-17
C_x_PM_AND3_X2__A1_c2 VSS N_A1_M0_g 7.76e-17
C_x_PM_AND3_X2__A1_c3 VSS N_A1_M4_g 4.58756e-17
R_x_PM_AND3_X2__A1_r4 x_PM_AND3_X2__A1_18 x_PM_AND3_X2__A1_14 4.74714
R_x_PM_AND3_X2__A1_r5 x_PM_AND3_X2__A1_17 x_PM_AND3_X2__A1_14 4.74714
R_x_PM_AND3_X2__A1_r6 x_PM_AND3_X2__A1_14 x_PM_AND3_X2__A1_12 25.0012
R_x_PM_AND3_X2__A1_r7 x_PM_AND3_X2__A1_12 A1 0.156071
R_x_PM_AND3_X2__A1_r8 N_A1_M0_g x_PM_AND3_X2__A1_18 106.47
R_x_PM_AND3_X2__A1_r9 N_A1_M4_g x_PM_AND3_X2__A1_17 42.9
C_x_PM_AND3_X2__A2_c0 VSS x_PM_AND3_X2__A2_14 8.59743e-18
C_x_PM_AND3_X2__A2_c1 VSS x_PM_AND3_X2__A2_12 5.83497e-17
C_x_PM_AND3_X2__A2_c2 VSS N_A2_M1_g 8.11148e-17
C_x_PM_AND3_X2__A2_c3 VSS N_A2_M5_g 4.54734e-17
R_x_PM_AND3_X2__A2_r4 x_PM_AND3_X2__A2_18 x_PM_AND3_X2__A2_14 4.7687
R_x_PM_AND3_X2__A2_r5 x_PM_AND3_X2__A2_17 x_PM_AND3_X2__A2_14 4.7687
R_x_PM_AND3_X2__A2_r6 x_PM_AND3_X2__A2_14 x_PM_AND3_X2__A2_12 25.0012
R_x_PM_AND3_X2__A2_r7 x_PM_AND3_X2__A2_12 A2 0.169643
R_x_PM_AND3_X2__A2_r8 N_A2_M1_g x_PM_AND3_X2__A2_18 106.47
R_x_PM_AND3_X2__A2_r9 N_A2_M5_g x_PM_AND3_X2__A2_17 42.9
C_x_PM_AND3_X2__A3_c0 VSS x_PM_AND3_X2__A3_14 8.46766e-18
C_x_PM_AND3_X2__A3_c1 VSS x_PM_AND3_X2__A3_12 5.10428e-17
C_x_PM_AND3_X2__A3_c2 VSS N_A3_M2_g 5.76331e-17
C_x_PM_AND3_X2__A3_c3 VSS N_A3_M6_g 6.8921e-17
R_x_PM_AND3_X2__A3_r4 x_PM_AND3_X2__A3_18 x_PM_AND3_X2__A3_14 4.7687
R_x_PM_AND3_X2__A3_r5 x_PM_AND3_X2__A3_17 x_PM_AND3_X2__A3_14 4.7687
R_x_PM_AND3_X2__A3_r6 x_PM_AND3_X2__A3_14 x_PM_AND3_X2__A3_12 25.0012
R_x_PM_AND3_X2__A3_r7 x_PM_AND3_X2__A3_12 A3 0.246296
R_x_PM_AND3_X2__A3_r8 N_A3_M2_g x_PM_AND3_X2__A3_18 67.47
R_x_PM_AND3_X2__A3_r9 N_A3_M6_g x_PM_AND3_X2__A3_17 81.9
C_x_PM_AND3_X2__ZN_c0 VSS N_ZN_M7_d 3.25194e-17
C_x_PM_AND3_X2__ZN_c1 VSS ZN 9.50381e-17
C_x_PM_AND3_X2__ZN_c2 VSS N_ZN_M3_d 5.591e-17
C_x_PM_AND3_X2__ZN_c3 VSS x_PM_AND3_X2__ZN_3 8.95839e-18
R_x_PM_AND3_X2__ZN_r4 ZN x_PM_AND3_X2__ZN_8 1.87286
R_x_PM_AND3_X2__ZN_r5 x_PM_AND3_X2__ZN_7 N_ZN_M7_d 0.30478
R_x_PM_AND3_X2__ZN_r6 ZN x_PM_AND3_X2__ZN_7 1.79143
R_x_PM_AND3_X2__ZN_r7 x_PM_AND3_X2__ZN_8 x_PM_AND3_X2__ZN_3 0.20978
R_x_PM_AND3_X2__ZN_r8 N_ZN_M3_d x_PM_AND3_X2__ZN_3 0.686111
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
