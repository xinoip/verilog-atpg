.SUBCKT and9 A1 A2 A3 A4 A5 A6 A7 A8 A9 VDD VSS ZN
**************************************************NAND3_X2***********************************************
M_M3 N_Zalp1_M0_d N_A3_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.037800P PS=0.750000U PD=0.820000U
M_M4 N_VDD_M1_d N_A2_M1_g N_Zalp1_M0_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.037800P PS=0.820000U PD=0.820000U
M_M5 N_Zalp1_M2_d N_A1_M2_g N_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 7 N_A3_M3_g N_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.340000U AS=0.035700P AD=0.047600P PS=0.890000U PD=0.960000U
M_M1 8 N_A2_M4_g 7 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.047600P PS=0.960000U PD=0.960000U
M_M2 N_Zalp1_M5_d N_A1_M5_g 8 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.035700P PS=0.960000U PD=0.890000U
C_x_PM_NAND3_X2__VSS_c0 VSS VSS 7.02872e-17
C_x_PM_NAND3_X2__VSS_c1 VSS x_PM_NAND3_X2__VSS_6 1.05487e-17
C_x_PM_NAND3_X2__VSS_c2 VSS N_VSS_M3_s 1.8134e-17
R_x_PM_NAND3_X2__VSS_r3 VSS x_PM_NAND3_X2__VSS_6 0.603529
R_x_PM_NAND3_X2__VSS_r4 x_PM_NAND3_X2__VSS_6 x_PM_NAND3_X2__VSS_2 0.264221
R_x_PM_NAND3_X2__VSS_r5 N_VSS_M3_s x_PM_NAND3_X2__VSS_2 0.230714
C_x_PM_NAND3_X2__VDD_c0 VSS N_VDD_M1_d 6.12848e-17
C_x_PM_NAND3_X2__VDD_c1 VSS x_PM_NAND3_X2__VDD_7 3.00804e-17
C_x_PM_NAND3_X2__VDD_c2 VSS N_VDD_M0_s 2.5125e-17
C_x_PM_NAND3_X2__VDD_c3 VSS x_PM_NAND3_X2__VDD_3 1.06055e-17
R_x_PM_NAND3_X2__VDD_r4 VDD x_PM_NAND3_X2__VDD_8 0.195294
R_x_PM_NAND3_X2__VDD_r5 x_PM_NAND3_X2__VDD_7 N_VDD_M1_d 0.140674
R_x_PM_NAND3_X2__VDD_r6 x_PM_NAND3_X2__VDD_8 x_PM_NAND3_X2__VDD_7 0.614706
R_x_PM_NAND3_X2__VDD_r7 VDD x_PM_NAND3_X2__VDD_3 0.0689273
R_x_PM_NAND3_X2__VDD_r8 N_VDD_M0_s x_PM_NAND3_X2__VDD_3 0.230714
C_x_PM_NAND3_X2__A3_c0 VSS x_PM_NAND3_X2__A3_14 6.68331e-18
C_x_PM_NAND3_X2__A3_c1 VSS x_PM_NAND3_X2__A3_12 3.18495e-17
C_x_PM_NAND3_X2__A3_c2 VSS N_A3_M0_g 7.81987e-17
C_x_PM_NAND3_X2__A3_c3 VSS N_A3_M3_g 4.14029e-17
R_x_PM_NAND3_X2__A3_r4 x_PM_NAND3_X2__A3_18 x_PM_NAND3_X2__A3_14 4.7687
R_x_PM_NAND3_X2__A3_r5 x_PM_NAND3_X2__A3_17 x_PM_NAND3_X2__A3_14 4.7687
R_x_PM_NAND3_X2__A3_r6 x_PM_NAND3_X2__A3_14 x_PM_NAND3_X2__A3_12 25.0012
R_x_PM_NAND3_X2__A3_r7 x_PM_NAND3_X2__A3_12 A3 0.0781486
R_x_PM_NAND3_X2__A3_r8 N_A3_M0_g x_PM_NAND3_X2__A3_18 95.94
R_x_PM_NAND3_X2__A3_r9 N_A3_M3_g x_PM_NAND3_X2__A3_17 35.1
C_x_PM_NAND3_X2__Zalp1_c0 VSS N_Zalp1_M5_d 1.32739e-16
C_x_PM_NAND3_X2__Zalp1_c1 VSS x_PM_NAND3_X2__Zalp1_8 1.01878e-17
C_x_PM_NAND3_X2__Zalp1_c2 VSS x_PM_NAND3_X2__Zalp1_4 7.15422e-17
R_x_PM_NAND3_X2__Zalp1_r3 Zalp1 N_Zalp1_M5_d 1.59389
R_x_PM_NAND3_X2__Zalp1_r4 N_Zalp1_M2_d x_PM_NAND3_X2__Zalp1_8 0.0406238
R_x_PM_NAND3_X2__Zalp1_r5 Zalp1 x_PM_NAND3_X2__Zalp1_8 1.28778
R_x_PM_NAND3_X2__Zalp1_r6 N_Zalp1_M2_d x_PM_NAND3_X2__Zalp1_4 0.176037
R_x_PM_NAND3_X2__Zalp1_r7 N_Zalp1_M0_d x_PM_NAND3_X2__Zalp1_4 1.85929
C_x_PM_NAND3_X2__A2_c0 VSS x_PM_NAND3_X2__A2_14 8.63262e-18
C_x_PM_NAND3_X2__A2_c1 VSS x_PM_NAND3_X2__A2_12 3.91329e-17
C_x_PM_NAND3_X2__A2_c2 VSS N_A2_M1_g 4.24405e-17
C_x_PM_NAND3_X2__A2_c3 VSS N_A2_M4_g 8.48173e-17
R_x_PM_NAND3_X2__A2_r4 x_PM_NAND3_X2__A2_18 x_PM_NAND3_X2__A2_14 4.7687
R_x_PM_NAND3_X2__A2_r5 x_PM_NAND3_X2__A2_17 x_PM_NAND3_X2__A2_14 4.7687
R_x_PM_NAND3_X2__A2_r6 x_PM_NAND3_X2__A2_14 x_PM_NAND3_X2__A2_12 25.0012
R_x_PM_NAND3_X2__A2_r7 x_PM_NAND3_X2__A2_12 A2 0.169643
R_x_PM_NAND3_X2__A2_r8 N_A2_M1_g x_PM_NAND3_X2__A2_18 29.64
R_x_PM_NAND3_X2__A2_r9 N_A2_M4_g x_PM_NAND3_X2__A2_17 101.4
C_x_PM_NAND3_X2__A1_c0 VSS x_PM_NAND3_X2__A1_18 1.22048e-17
C_x_PM_NAND3_X2__A1_c1 VSS x_PM_NAND3_X2__A1_12 7.61168e-17
C_x_PM_NAND3_X2__A1_c2 VSS N_A1_M2_g 8.98944e-17
C_x_PM_NAND3_X2__A1_c3 VSS N_A1_M5_g 4.86035e-17
R_x_PM_NAND3_X2__A1_r4 x_PM_NAND3_X2__A1_18 x_PM_NAND3_X2__A1_14 3.9
R_x_PM_NAND3_X2__A1_r5 x_PM_NAND3_X2__A1_14 x_PM_NAND3_X2__A1_12 25.0012
R_x_PM_NAND3_X2__A1_r6 x_PM_NAND3_X2__A1_12 A1 0.0459677
R_x_PM_NAND3_X2__A1_r7 x_PM_NAND3_X2__A1_18 x_PM_NAND3_X2__A1_5 1.95
R_x_PM_NAND3_X2__A1_r8 N_A1_M2_g x_PM_NAND3_X2__A1_5 95.94
R_x_PM_NAND3_X2__A1_r9 x_PM_NAND3_X2__A1_18 x_PM_NAND3_X2__A1_VSS 1.95
R_x_PM_NAND3_X2__A1_r10 N_A1_M5_g x_PM_NAND3_X2__A1_VSS 35.1

**************************************************NAND3_X2***********************************************
M2_M3 N2_Zalp2_M0_d N2_A6_M0_g N2_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.037800P PS=0.750000U PD=0.820000U
M2_M4 N2_VDD_M1_d N2_A5_M1_g N2_Zalp2_M0_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.037800P PS=0.820000U PD=0.820000U
M2_M5 N2_Zalp2_M2_d N2_A4_M2_g N2_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.028350P PS=0.820000U PD=0.750000U
M2_M0 72 N2_A6_M3_g N2_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.340000U AS=0.035700P AD=0.047600P PS=0.890000U PD=0.960000U
M2_M1 82 N2_A5_M4_g 72 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.047600P PS=0.960000U PD=0.960000U
M2_M2 N2_Zalp2_M5_d N2_A4_M5_g 82 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.035700P PS=0.960000U PD=0.890000U
C_x2_PM2_NAND3_X2__VSS_c0 VSS VSS 7.02872e-17
C_x2_PM2_NAND3_X2__VSS_c1 VSS x2_PM2_NAND3_X2__VSS_6 1.05487e-17
C_x2_PM2_NAND3_X2__VSS_c2 VSS N2_VSS_M3_s 1.8134e-17
R_x2_PM2_NAND3_X2__VSS_r3 VSS x2_PM2_NAND3_X2__VSS_6 0.603529
R_x2_PM2_NAND3_X2__VSS_r4 x2_PM2_NAND3_X2__VSS_6 x2_PM2_NAND3_X2__VSS_2 0.264221
R_x2_PM2_NAND3_X2__VSS_r5 N2_VSS_M3_s x2_PM2_NAND3_X2__VSS_2 0.230714
C_x2_PM2_NAND3_X2__VDD_c0 VSS N2_VDD_M1_d 6.12848e-17
C_x2_PM2_NAND3_X2__VDD_c1 VSS x2_PM2_NAND3_X2__VDD_7 3.00804e-17
C_x2_PM2_NAND3_X2__VDD_c2 VSS N2_VDD_M0_s 2.5125e-17
C_x2_PM2_NAND3_X2__VDD_c3 VSS x2_PM2_NAND3_X2__VDD_3 1.06055e-17
R_x2_PM2_NAND3_X2__VDD_r4 VDD x2_PM2_NAND3_X2__VDD_8 0.195294
R_x2_PM2_NAND3_X2__VDD_r5 x2_PM2_NAND3_X2__VDD_7 N2_VDD_M1_d 0.140674
R_x2_PM2_NAND3_X2__VDD_r6 x2_PM2_NAND3_X2__VDD_8 x2_PM2_NAND3_X2__VDD_7 0.614706
R_x2_PM2_NAND3_X2__VDD_r7 VDD x2_PM2_NAND3_X2__VDD_3 0.0689273
R_x2_PM2_NAND3_X2__VDD_r8 N2_VDD_M0_s x2_PM2_NAND3_X2__VDD_3 0.230714
C_x2_PM2_NAND3_X2__A6_c0 VSS x2_PM2_NAND3_X2__A6_14 6.68331e-18
C_x2_PM2_NAND3_X2__A6_c1 VSS x2_PM2_NAND3_X2__A6_12 3.18495e-17
C_x2_PM2_NAND3_X2__A6_c2 VSS N2_A6_M0_g 7.81987e-17
C_x2_PM2_NAND3_X2__A6_c3 VSS N2_A6_M3_g 4.14029e-17
R_x2_PM2_NAND3_X2__A6_r4 x2_PM2_NAND3_X2__A6_18 x2_PM2_NAND3_X2__A6_14 4.7687
R_x2_PM2_NAND3_X2__A6_r5 x2_PM2_NAND3_X2__A6_17 x2_PM2_NAND3_X2__A6_14 4.7687
R_x2_PM2_NAND3_X2__A6_r6 x2_PM2_NAND3_X2__A6_14 x2_PM2_NAND3_X2__A6_12 25.0012
R_x2_PM2_NAND3_X2__A6_r7 x2_PM2_NAND3_X2__A6_12 A6 0.0781486
R_x2_PM2_NAND3_X2__A6_r8 N2_A6_M0_g x2_PM2_NAND3_X2__A6_18 95.94
R_x2_PM2_NAND3_X2__A6_r9 N2_A6_M3_g x2_PM2_NAND3_X2__A6_17 35.1
C_x2_PM2_NAND3_X2__Zalp2_c0 VSS N2_Zalp2_M5_d 1.32739e-16
C_x2_PM2_NAND3_X2__Zalp2_c1 VSS x2_PM2_NAND3_X2__Zalp2_8 1.01878e-17
C_x2_PM2_NAND3_X2__Zalp2_c2 VSS x2_PM2_NAND3_X2__Zalp2_4 7.15422e-17
R_x2_PM2_NAND3_X2__Zalp2_r3 Zalp2 N2_Zalp2_M5_d 1.59389
R_x2_PM2_NAND3_X2__Zalp2_r4 N2_Zalp2_M2_d x2_PM2_NAND3_X2__Zalp2_8 0.0406238
R_x2_PM2_NAND3_X2__Zalp2_r5 Zalp2 x2_PM2_NAND3_X2__Zalp2_8 1.28778
R_x2_PM2_NAND3_X2__Zalp2_r6 N2_Zalp2_M2_d x2_PM2_NAND3_X2__Zalp2_4 0.176037
R_x2_PM2_NAND3_X2__Zalp2_r7 N2_Zalp2_M0_d x2_PM2_NAND3_X2__Zalp2_4 1.85929
C_x2_PM2_NAND3_X2__A5_c0 VSS x2_PM2_NAND3_X2__A5_14 8.63262e-18
C_x2_PM2_NAND3_X2__A5_c1 VSS x2_PM2_NAND3_X2__A5_12 3.91329e-17
C_x2_PM2_NAND3_X2__A5_c2 VSS N2_A5_M1_g 4.24405e-17
C_x2_PM2_NAND3_X2__A5_c3 VSS N2_A5_M4_g 8.48173e-17
R_x2_PM2_NAND3_X2__A5_r4 x2_PM2_NAND3_X2__A5_18 x2_PM2_NAND3_X2__A5_14 4.7687
R_x2_PM2_NAND3_X2__A5_r5 x2_PM2_NAND3_X2__A5_17 x2_PM2_NAND3_X2__A5_14 4.7687
R_x2_PM2_NAND3_X2__A5_r6 x2_PM2_NAND3_X2__A5_14 x2_PM2_NAND3_X2__A5_12 25.0012
R_x2_PM2_NAND3_X2__A5_r7 x2_PM2_NAND3_X2__A5_12 A5 0.169643
R_x2_PM2_NAND3_X2__A5_r8 N2_A5_M1_g x2_PM2_NAND3_X2__A5_18 29.64
R_x2_PM2_NAND3_X2__A5_r9 N2_A5_M4_g x2_PM2_NAND3_X2__A5_17 101.4
C_x2_PM2_NAND3_X2__A4_c0 VSS x2_PM2_NAND3_X2__A4_18 1.22048e-17
C_x2_PM2_NAND3_X2__A4_c1 VSS x2_PM2_NAND3_X2__A4_12 7.61168e-17
C_x2_PM2_NAND3_X2__A4_c2 VSS N2_A4_M2_g 8.98944e-17
C_x2_PM2_NAND3_X2__A4_c3 VSS N2_A4_M5_g 4.86035e-17
R_x2_PM2_NAND3_X2__A4_r4 x2_PM2_NAND3_X2__A4_18 x2_PM2_NAND3_X2__A4_14 3.9
R_x2_PM2_NAND3_X2__A4_r5 x2_PM2_NAND3_X2__A4_14 x2_PM2_NAND3_X2__A4_12 25.0012
R_x2_PM2_NAND3_X2__A4_r6 x2_PM2_NAND3_X2__A4_12 A4 0.0459677
R_x2_PM2_NAND3_X2__A4_r7 x2_PM2_NAND3_X2__A4_18 x2_PM2_NAND3_X2__A4_5 1.95
R_x2_PM2_NAND3_X2__A4_r8 N2_A4_M2_g x2_PM2_NAND3_X2__A4_5 95.94
R_x2_PM2_NAND3_X2__A4_r9 x2_PM2_NAND3_X2__A4_18 x2_PM2_NAND3_X2__A4_VSS 1.95
R_x2_PM2_NAND3_X2__A4_r10 N2_A4_M5_g x2_PM2_NAND3_X2__A4_VSS 35.1

**************************************************NAND3_X2***********************************************
M3_M3 N3_Zalp3_M0_d N3_A9_M0_g N3_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.037800P PS=0.750000U PD=0.820000U
M3_M4 N3_VDD_M1_d N3_A8_M1_g N3_Zalp3_M0_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.037800P PS=0.820000U PD=0.820000U
M3_M5 N3_Zalp3_M2_d N3_A7_M2_g N3_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.028350P PS=0.820000U PD=0.750000U
M3_M0 73 N3_A9_M3_g N3_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.340000U AS=0.035700P AD=0.047600P PS=0.890000U PD=0.960000U
M3_M1 83 N3_A8_M4_g 73 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.047600P PS=0.960000U PD=0.960000U
M3_M2 N3_Zalp3_M5_d N3_A7_M5_g 83 VSS NMOS_VTL L=0.050U W=0.340000U AS=0.047600P AD=0.035700P PS=0.960000U PD=0.890000U
C_x3_PM3_NAND3_X2__VSS_c0 VSS VSS 7.02872e-17
C_x3_PM3_NAND3_X2__VSS_c1 VSS x3_PM3_NAND3_X2__VSS_6 1.05487e-17
C_x3_PM3_NAND3_X2__VSS_c2 VSS N3_VSS_M3_s 1.8134e-17
R_x3_PM3_NAND3_X2__VSS_r3 VSS x3_PM3_NAND3_X2__VSS_6 0.603529
R_x3_PM3_NAND3_X2__VSS_r4 x3_PM3_NAND3_X2__VSS_6 x3_PM3_NAND3_X2__VSS_2 0.264221
R_x3_PM3_NAND3_X2__VSS_r5 N3_VSS_M3_s x3_PM3_NAND3_X2__VSS_2 0.230714
C_x3_PM3_NAND3_X2__VDD_c0 VSS N3_VDD_M1_d 6.12848e-17
C_x3_PM3_NAND3_X2__VDD_c1 VSS x3_PM3_NAND3_X2__VDD_7 3.00804e-17
C_x3_PM3_NAND3_X2__VDD_c2 VSS N3_VDD_M0_s 2.5125e-17
C_x3_PM3_NAND3_X2__VDD_c3 VSS x3_PM3_NAND3_X2__VDD_3 1.06055e-17
R_x3_PM3_NAND3_X2__VDD_r4 VDD x3_PM3_NAND3_X2__VDD_8 0.195294
R_x3_PM3_NAND3_X2__VDD_r5 x3_PM3_NAND3_X2__VDD_7 N3_VDD_M1_d 0.140674
R_x3_PM3_NAND3_X2__VDD_r6 x3_PM3_NAND3_X2__VDD_8 x3_PM3_NAND3_X2__VDD_7 0.614706
R_x3_PM3_NAND3_X2__VDD_r7 VDD x3_PM3_NAND3_X2__VDD_3 0.0689273
R_x3_PM3_NAND3_X2__VDD_r8 N3_VDD_M0_s x3_PM3_NAND3_X2__VDD_3 0.230714
C_x3_PM3_NAND3_X2__A9_c0 VSS x3_PM3_NAND3_X2__A9_14 6.68331e-18
C_x3_PM3_NAND3_X2__A9_c1 VSS x3_PM3_NAND3_X2__A9_12 3.18495e-17
C_x3_PM3_NAND3_X2__A9_c2 VSS N3_A9_M0_g 7.81987e-17
C_x3_PM3_NAND3_X2__A9_c3 VSS N3_A9_M3_g 4.14029e-17
R_x3_PM3_NAND3_X2__A9_r4 x3_PM3_NAND3_X2__A9_18 x3_PM3_NAND3_X2__A9_14 4.7687
R_x3_PM3_NAND3_X2__A9_r5 x3_PM3_NAND3_X2__A9_17 x3_PM3_NAND3_X2__A9_14 4.7687
R_x3_PM3_NAND3_X2__A9_r6 x3_PM3_NAND3_X2__A9_14 x3_PM3_NAND3_X2__A9_12 25.0012
R_x3_PM3_NAND3_X2__A9_r7 x3_PM3_NAND3_X2__A9_12 A9 0.0781486
R_x3_PM3_NAND3_X2__A9_r8 N3_A9_M0_g x3_PM3_NAND3_X2__A9_18 95.94
R_x3_PM3_NAND3_X2__A9_r9 N3_A9_M3_g x3_PM3_NAND3_X2__A9_17 35.1
C_x3_PM3_NAND3_X2__Zalp3_c0 VSS N3_Zalp3_M5_d 1.32739e-16
C_x3_PM3_NAND3_X2__Zalp3_c1 VSS x3_PM3_NAND3_X2__Zalp3_8 1.01878e-17
C_x3_PM3_NAND3_X2__Zalp3_c2 VSS x3_PM3_NAND3_X2__Zalp3_4 7.15422e-17
R_x3_PM3_NAND3_X2__Zalp3_r3 Zalp3 N3_Zalp3_M5_d 1.59389
R_x3_PM3_NAND3_X2__Zalp3_r4 N3_Zalp3_M2_d x3_PM3_NAND3_X2__Zalp3_8 0.0406238
R_x3_PM3_NAND3_X2__Zalp3_r5 Zalp3 x3_PM3_NAND3_X2__Zalp3_8 1.28778
R_x3_PM3_NAND3_X2__Zalp3_r6 N3_Zalp3_M2_d x3_PM3_NAND3_X2__Zalp3_4 0.176037
R_x3_PM3_NAND3_X2__Zalp3_r7 N3_Zalp3_M0_d x3_PM3_NAND3_X2__Zalp3_4 1.85929
C_x3_PM3_NAND3_X2__A8_c0 VSS x3_PM3_NAND3_X2__A8_14 8.63262e-18
C_x3_PM3_NAND3_X2__A8_c1 VSS x3_PM3_NAND3_X2__A8_12 3.91329e-17
C_x3_PM3_NAND3_X2__A8_c2 VSS N3_A8_M1_g 4.24405e-17
C_x3_PM3_NAND3_X2__A8_c3 VSS N3_A8_M4_g 8.48173e-17
R_x3_PM3_NAND3_X2__A8_r4 x3_PM3_NAND3_X2__A8_18 x3_PM3_NAND3_X2__A8_14 4.7687
R_x3_PM3_NAND3_X2__A8_r5 x3_PM3_NAND3_X2__A8_17 x3_PM3_NAND3_X2__A8_14 4.7687
R_x3_PM3_NAND3_X2__A8_r6 x3_PM3_NAND3_X2__A8_14 x3_PM3_NAND3_X2__A8_12 25.0012
R_x3_PM3_NAND3_X2__A8_r7 x3_PM3_NAND3_X2__A8_12 A8 0.169643
R_x3_PM3_NAND3_X2__A8_r8 N3_A8_M1_g x3_PM3_NAND3_X2__A8_18 29.64
R_x3_PM3_NAND3_X2__A8_r9 N3_A8_M4_g x3_PM3_NAND3_X2__A8_17 101.4
C_x3_PM3_NAND3_X2__A7_c0 VSS x3_PM3_NAND3_X2__A7_18 1.22048e-17
C_x3_PM3_NAND3_X2__A7_c1 VSS x3_PM3_NAND3_X2__A7_12 7.61168e-17
C_x3_PM3_NAND3_X2__A7_c2 VSS N3_A7_M2_g 8.98944e-17
C_x3_PM3_NAND3_X2__A7_c3 VSS N3_A7_M5_g 4.86035e-17
R_x3_PM3_NAND3_X2__A7_r4 x3_PM3_NAND3_X2__A7_18 x3_PM3_NAND3_X2__A7_14 3.9
R_x3_PM3_NAND3_X2__A7_r5 x3_PM3_NAND3_X2__A7_14 x3_PM3_NAND3_X2__A7_12 25.0012
R_x3_PM3_NAND3_X2__A7_r6 x3_PM3_NAND3_X2__A7_12 A7 0.0459677
R_x3_PM3_NAND3_X2__A7_r7 x3_PM3_NAND3_X2__A7_18 x3_PM3_NAND3_X2__A7_5 1.95
R_x3_PM3_NAND3_X2__A7_r8 N3_A7_M2_g x3_PM3_NAND3_X2__A7_5 95.94
R_x3_PM3_NAND3_X2__A7_r9 x3_PM3_NAND3_X2__A7_18 x3_PM3_NAND3_X2__A7_VSS 1.95
R_x3_PM3_NAND3_X2__A7_r10 N3_A7_M5_g x3_PM3_NAND3_X2__A7_VSS 35.1

*********************************************NOR3_X2*************************************************************
M4_M3 74 N4_Zalp3_M0_g N4_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.520000U AS=0.054600P AD=0.072800P PS=1.250000U PD=1.320000U
M4_M4 84 N4_Zalp2_M1_g 74 VDD PMOS_VTL L=0.050U W=0.520000U AS=0.072800P AD=0.072800P PS=1.320000U PD=1.320000U
M4_M5 N4_ZN4_M2_d N4_Zalp1_M2_g 84 VDD PMOS_VTL L=0.050U W=0.520000U AS=0.072800P AD=0.054600P PS=1.320000U PD=1.250000U
M4_M0 N4_ZN4_M3_d N4_Zalp3_M3_g N4_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M4_M1 N4_VSS_M4_d N4_Zalp2_M4_g N4_ZN4_M3_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.025200P PS=0.640000U PD=0.640000U
M4_M2 N4_ZN4_M5_d N4_Zalp1_M5_g N4_VSS_M4_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x4_PM_NOR3_X2__VSS_c0 VSS x4_PM_NOR3_X2__VSS_17 4.46075e-17
C_x4_PM_NOR3_X2__VSS_c1 VSS N4_VSS_M4_d 2.78358e-17
C_x4_PM_NOR3_X2__VSS_c2 VSS x4_PM_NOR3_X2__VSS_8 1.05487e-17
C_x4_PM_NOR3_X2__VSS_c3 VSS x4_PM_NOR3_X2__VSS_7 3.86305e-17
C_x4_PM_NOR3_X2__VSS_c4 VSS N4_VSS_M3_s 9.87304e-18
R_x4_PM_NOR3_X2__VSS_r5 x4_PM_NOR3_X2__VSS_17 x4_PM_NOR3_X2__VSS_11 0.145286
R_x4_PM_NOR3_X2__VSS_r6 N4_VSS_M4_d x4_PM_NOR3_X2__VSS_11 0.230714
R_x4_PM_NOR3_X2__VSS_r7 VSS x4_PM_NOR3_X2__VSS_8 0.603529
R_x4_PM_NOR3_X2__VSS_r8 x4_PM_NOR3_X2__VSS_17 x4_PM_NOR3_X2__VSS_7 0.0731438
R_x4_PM_NOR3_X2__VSS_r9 VSS x4_PM_NOR3_X2__VSS_7 0.0782353
R_x4_PM_NOR3_X2__VSS_r10 x4_PM_NOR3_X2__VSS_8 x4_PM_NOR3_X2__VSS_3 0.264221
R_x4_PM_NOR3_X2__VSS_r11 N4_VSS_M3_s x4_PM_NOR3_X2__VSS_3 0.230714
C_x4_PM_NOR3_X2__VDD_c0 VSS VDD 5.9596e-17
C_x4_PM_NOR3_X2__VDD_c1 VSS N4_VDD_M0_s 2.58417e-17
C_x4_PM_NOR3_X2__VDD_c2 VSS x4_PM_NOR3_X2__VDD_2 1.06055e-17
R_x4_PM_NOR3_X2__VDD_r3 VDD x4_PM_NOR3_X2__VDD_2 0.0689273
R_x4_PM_NOR3_X2__VDD_r4 N4_VDD_M0_s x4_PM_NOR3_X2__VDD_2 0.230714
C_x4_PM_NOR3_X2__Zalp3_c0 VSS x4_PM_NOR3_X2__Zalp3_11 7.14715e-18
C_x4_PM_NOR3_X2__Zalp3_c1 VSS x4_PM_NOR3_X2__Zalp3_9 5.04542e-17
C_x4_PM_NOR3_X2__Zalp3_c2 VSS N4_Zalp3_M0_g 6.20936e-17
C_x4_PM_NOR3_X2__Zalp3_c3 VSS N4_Zalp3_M3_g 5.91756e-17
R_x4_PM_NOR3_X2__Zalp3_r4 x4_PM_NOR3_X2__Zalp3_18 x4_PM_NOR3_X2__Zalp3_11 4.74714
R_x4_PM_NOR3_X2__Zalp3_r5 x4_PM_NOR3_X2__Zalp3_17 x4_PM_NOR3_X2__Zalp3_11 4.74714
R_x4_PM_NOR3_X2__Zalp3_r6 x4_PM_NOR3_X2__Zalp3_11 x4_PM_NOR3_X2__Zalp3_9 25.0012
R_x4_PM_NOR3_X2__Zalp3_r7 Zalp3 x4_PM_NOR3_X2__Zalp3_9 0.2204
R_x4_PM_NOR3_X2__Zalp3_r8 N4_Zalp3_M0_g x4_PM_NOR3_X2__Zalp3_18 49.14
R_x4_PM_NOR3_X2__Zalp3_r9 N4_Zalp3_M3_g x4_PM_NOR3_X2__Zalp3_17 74.88
C_x4_PM_NOR3_X2__ZN4_c0 VSS x4_PM_NOR3_X2__ZN4_22 2.56413e-18
C_x4_PM_NOR3_X2__ZN4_c1 VSS ZN 5.06951e-17
C_x4_PM_NOR3_X2__ZN4_c2 VSS N4_ZN4_M2_d 2.75881e-17
C_x4_PM_NOR3_X2__ZN4_c3 VSS x4_PM_NOR3_X2__ZN4_14 6.25994e-18
C_x4_PM_NOR3_X2__ZN4_c4 VSS N4_ZN4_M5_d 2.52851e-17
C_x4_PM_NOR3_X2__ZN4_c5 VSS x4_PM_NOR3_X2__ZN4_9 8.16416e-18
C_x4_PM_NOR3_X2__ZN4_c6 VSS x4_PM_NOR3_X2__ZN4_8 4.12951e-17
C_x4_PM_NOR3_X2__ZN4_c7 VSS N4_ZN4_M3_d 2.15312e-17
R_x4_PM_NOR3_X2__ZN4_r8 ZN x4_PM_NOR3_X2__ZN4_19 1.46571
R_x4_PM_NOR3_X2__ZN4_r9 x4_PM_NOR3_X2__ZN4_22 x4_PM_NOR3_X2__ZN4_18 0.143785
R_x4_PM_NOR3_X2__ZN4_r10 ZN x4_PM_NOR3_X2__ZN4_18 0.868571
R_x4_PM_NOR3_X2__ZN4_r11 x4_PM_NOR3_X2__ZN4_19 x4_PM_NOR3_X2__ZN4_14 0.20978
R_x4_PM_NOR3_X2__ZN4_r12 N4_ZN4_M2_d x4_PM_NOR3_X2__ZN4_14 0.686111
R_x4_PM_NOR3_X2__ZN4_r13 x4_PM_NOR3_X2__ZN4_22 x4_PM_NOR3_X2__ZN4_10 0.143785
R_x4_PM_NOR3_X2__ZN4_r14 N4_ZN4_M5_d x4_PM_NOR3_X2__ZN4_10 0.116111
R_x4_PM_NOR3_X2__ZN4_r15 x4_PM_NOR3_X2__ZN4_22 x4_PM_NOR3_X2__ZN4_8 0.0569232
R_x4_PM_NOR3_X2__ZN4_r16 x4_PM_NOR3_X2__ZN4_9 x4_PM_NOR3_X2__ZN4_8 1.65571
R_x4_PM_NOR3_X2__ZN4_r17 x4_PM_NOR3_X2__ZN4_9 x4_PM_NOR3_X2__ZN4_4 0.212317
R_x4_PM_NOR3_X2__ZN4_r18 N4_ZN4_M3_d x4_PM_NOR3_X2__ZN4_4 0.149286
C_x4_PM_NOR3_X2__Zalp2_c0 VSS x4_PM_NOR3_X2__Zalp2_11 8.98632e-18
C_x4_PM_NOR3_X2__Zalp2_c1 VSS x4_PM_NOR3_X2__Zalp2_9 8.53584e-17
C_x4_PM_NOR3_X2__Zalp2_c2 VSS N4_Zalp2_M1_g 6.12109e-17
C_x4_PM_NOR3_X2__Zalp2_c3 VSS N4_Zalp2_M4_g 6.60015e-17
R_x4_PM_NOR3_X2__Zalp2_r4 x4_PM_NOR3_X2__Zalp2_18 x4_PM_NOR3_X2__Zalp2_11 4.74714
R_x4_PM_NOR3_X2__Zalp2_r5 x4_PM_NOR3_X2__Zalp2_17 x4_PM_NOR3_X2__Zalp2_11 4.74714
R_x4_PM_NOR3_X2__Zalp2_r6 x4_PM_NOR3_X2__Zalp2_11 x4_PM_NOR3_X2__Zalp2_9 25.0012
R_x4_PM_NOR3_X2__Zalp2_r7 Zalp2 x4_PM_NOR3_X2__Zalp2_9 0.2204
R_x4_PM_NOR3_X2__Zalp2_r8 N4_Zalp2_M1_g x4_PM_NOR3_X2__Zalp2_18 49.14
R_x4_PM_NOR3_X2__Zalp2_r9 N4_Zalp2_M4_g x4_PM_NOR3_X2__Zalp2_17 74.88
C_x4_PM_NOR3_X2__Zalp1_c0 VSS x4_PM_NOR3_X2__Zalp1_20 1.07269e-17
C_x4_PM_NOR3_X2__Zalp1_c1 VSS x4_PM_NOR3_X2__Zalp1_14 4.59258e-17
C_x4_PM_NOR3_X2__Zalp1_c2 VSS x4_PM_NOR3_X2__Zalp1_9 3.45973e-17
C_x4_PM_NOR3_X2__Zalp1_c3 VSS N4_Zalp1_M2_g 7.00434e-17
C_x4_PM_NOR3_X2__Zalp1_c4 VSS N4_Zalp1_M5_g 6.63408e-17
R_x4_PM_NOR3_X2__Zalp1_r5 x4_PM_NOR3_X2__Zalp1_20 x4_PM_NOR3_X2__Zalp1_16 2.34
R_x4_PM_NOR3_X2__Zalp1_r6 x4_PM_NOR3_X2__Zalp1_16 x4_PM_NOR3_X2__Zalp1_14 25.0012
R_x4_PM_NOR3_X2__Zalp1_r7 x4_PM_NOR3_X2__Zalp1_14 x4_PM_NOR3_X2__Zalp1_12 0.147778
R_x4_PM_NOR3_X2__Zalp1_r8 x4_PM_NOR3_X2__Zalp1_12 x4_PM_NOR3_X2__Zalp1_9 0.095
R_x4_PM_NOR3_X2__Zalp1_r9 Zalp1 x4_PM_NOR3_X2__Zalp1_9 0.298571
R_x4_PM_NOR3_X2__Zalp1_r10 x4_PM_NOR3_X2__Zalp1_20 x4_PM_NOR3_X2__Zalp1_5 1.95
R_x4_PM_NOR3_X2__Zalp1_r11 N4_Zalp1_M2_g x4_PM_NOR3_X2__Zalp1_5 56.94
R_x4_PM_NOR3_X2__Zalp1_r12 x4_PM_NOR3_X2__Zalp1_20 x4_PM_NOR3_X2__Zalp1_VSS 1.95
R_x4_PM_NOR3_X2__Zalp1_r13 N4_Zalp1_M5_g x4_PM_NOR3_X2__Zalp1_VSS 67.08
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
