.SUBCKT nor2 A1 A2 VDD VSS ZN  
M_M2 6 N_A2_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.390000U AS=0.040950P AD=0.054600P PS=0.990000U PD=1.060000U
M_M3 N_ZN_M1_d N_A1_M1_g 6 VDD PMOS_VTL L=0.050U W=0.390000U AS=0.054600P AD=0.040950P PS=1.060000U PD=0.990000U
M_M0 N_ZN_M2_d N_A2_M2_g N_VSS_M2_s VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.025200P PS=0.570000U PD=0.640000U
M_M1 N_VSS_M3_d N_A1_M3_g N_ZN_M2_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.025200P AD=0.018900P PS=0.640000U PD=0.570000U
C_x_PM_NOR2_X2__VSS_c0 VSS N_VSS_M3_d 1.9003e-17
C_x_PM_NOR2_X2__VSS_c1 VSS x_PM_NOR2_X2__VSS_8 1.14613e-17
C_x_PM_NOR2_X2__VSS_c2 VSS x_PM_NOR2_X2__VSS_7 5.12113e-17
C_x_PM_NOR2_X2__VSS_c3 VSS N_VSS_M2_s 1.7976e-17
R_x_PM_NOR2_X2__VSS_r4 N_VSS_M3_d x_PM_NOR2_X2__VSS_11 0.230714
R_x_PM_NOR2_X2__VSS_r5 VSS x_PM_NOR2_X2__VSS_8 0.357647
R_x_PM_NOR2_X2__VSS_r6 x_PM_NOR2_X2__VSS_11 x_PM_NOR2_X2__VSS_7 0.264221
R_x_PM_NOR2_X2__VSS_r7 VSS x_PM_NOR2_X2__VSS_7 0.324118
R_x_PM_NOR2_X2__VSS_r8 x_PM_NOR2_X2__VSS_8 x_PM_NOR2_X2__VSS_3 0.264221
R_x_PM_NOR2_X2__VSS_r9 N_VSS_M2_s x_PM_NOR2_X2__VSS_3 0.230714
C_x_PM_NOR2_X2__VDD_c0 VSS VDD 5.55967e-17
C_x_PM_NOR2_X2__VDD_c1 VSS N_VDD_M0_s 2.30938e-17
R_x_PM_NOR2_X2__VDD_r2 x_PM_NOR2_X2__VDD_10 VDD 0.0881799
R_x_PM_NOR2_X2__VDD_r3 N_VDD_M0_s x_PM_NOR2_X2__VDD_10 0.230714
C_x_PM_NOR2_X2__A2_c0 VSS x_PM_NOR2_X2__A2_18 8.24826e-18
C_x_PM_NOR2_X2__A2_c1 VSS x_PM_NOR2_X2__A2_12 4.45792e-17
C_x_PM_NOR2_X2__A2_c2 VSS N_A2_M0_g 9.21574e-17
C_x_PM_NOR2_X2__A2_c3 VSS N_A2_M2_g 3.09335e-17
R_x_PM_NOR2_X2__A2_r4 x_PM_NOR2_X2__A2_18 x_PM_NOR2_X2__A2_14 3.38
R_x_PM_NOR2_X2__A2_r5 x_PM_NOR2_X2__A2_14 x_PM_NOR2_X2__A2_12 25.0012
R_x_PM_NOR2_X2__A2_r6 x_PM_NOR2_X2__A2_12 A2 0.15069
R_x_PM_NOR2_X2__A2_r7 x_PM_NOR2_X2__A2_18 x_PM_NOR2_X2__A2_5 1.95
R_x_PM_NOR2_X2__A2_r8 N_A2_M0_g x_PM_NOR2_X2__A2_5 112.32
R_x_PM_NOR2_X2__A2_r9 x_PM_NOR2_X2__A2_18 x_PM_NOR2_X2__A2_VSS 1.95
R_x_PM_NOR2_X2__A2_r10 N_A2_M2_g x_PM_NOR2_X2__A2_VSS 21.84
C_x_PM_NOR2_X2__ZN_c0 VSS N_ZN_M1_d 5.96075e-17
C_x_PM_NOR2_X2__ZN_c1 VSS x_PM_NOR2_X2__ZN_9 3.74417e-17
C_x_PM_NOR2_X2__ZN_c2 VSS ZN 7.19517e-18
C_x_PM_NOR2_X2__ZN_c3 VSS N_ZN_M2_d 8.47483e-17
R_x_PM_NOR2_X2__ZN_r4 N_ZN_M1_d x_PM_NOR2_X2__ZN_11 2.91786
R_x_PM_NOR2_X2__ZN_r5 x_PM_NOR2_X2__ZN_11 x_PM_NOR2_X2__ZN_9 0.212317
R_x_PM_NOR2_X2__ZN_r6 x_PM_NOR2_X2__ZN_10 x_PM_NOR2_X2__ZN_9 0.597143
R_x_PM_NOR2_X2__ZN_r7 x_PM_NOR2_X2__ZN_10 ZN 0.212317
R_x_PM_NOR2_X2__ZN_r8 ZN x_PM_NOR2_X2__ZN_7 0.000542857
R_x_PM_NOR2_X2__ZN_r9 x_PM_NOR2_X2__ZN_7 N_ZN_M2_d 1.39731
C_x_PM_NOR2_X2__A1_c0 VSS A1 6.50458e-17
C_x_PM_NOR2_X2__A1_c1 VSS x_PM_NOR2_X2__A1_11 9.81933e-18
C_x_PM_NOR2_X2__A1_c2 VSS N_A1_M1_g 1.07185e-16
C_x_PM_NOR2_X2__A1_c3 VSS N_A1_M3_g 3.09279e-17
R_x_PM_NOR2_X2__A1_r4 x_PM_NOR2_X2__A1_11 x_PM_NOR2_X2__A1_16 4.42
R_x_PM_NOR2_X2__A1_r5 x_PM_NOR2_X2__A1_11 x_PM_NOR2_X2__A1_9 25.0012
R_x_PM_NOR2_X2__A1_r6 A1 x_PM_NOR2_X2__A1_9 0.15069
R_x_PM_NOR2_X2__A1_r7 x_PM_NOR2_X2__A1_16 x_PM_NOR2_X2__A1_5 1.95
R_x_PM_NOR2_X2__A1_r8 N_A1_M1_g x_PM_NOR2_X2__A1_5 112.32
R_x_PM_NOR2_X2__A1_r9 x_PM_NOR2_X2__A1_16 x_PM_NOR2_X2__A1_VSS 1.95
R_x_PM_NOR2_X2__A1_r10 N_A1_M3_g x_PM_NOR2_X2__A1_VSS 21.84
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
