.SUBCKT xor2 A B VDD VSS Z 
M_M5 8 N_A_M0_g N_3_M0_s VDD PMOS_VTL L=0.050U W=0.195000U AS=0.020475P AD=0.027300P PS=0.600000U PD=0.670000U
M_M6 N_VDD_M1_d N_B_M1_g 8 VDD PMOS_VTL L=0.050U W=0.195000U AS=0.027300P AD=0.040950P PS=0.670000U PD=1.060000U
M_M7 N_7_M2_d N_3_M2_g N_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.390000U AS=0.040950P AD=0.060450P PS=1.060000U PD=1.090000U
M_M8 N_Z_M3_d N_A_M3_g N_7_M2_d VDD PMOS_VTL L=0.050U W=0.390000U AS=0.060450P AD=0.054600P PS=1.090000U PD=1.060000U
M_M9 N_7_M4_d N_B_M4_g N_Z_M3_d VDD PMOS_VTL L=0.050U W=0.390000U AS=0.054600P AD=0.040950P PS=1.060000U PD=0.990000U
M_M0 N_3_M5_d N_A_M5_g N_VSS_M5_s VSS NMOS_VTL L=0.050U W=0.090000U AS=0.009450P AD=0.012600P PS=0.390000U PD=0.460000U
M_M1 N_VSS_M6_d N_B_M6_g N_3_M5_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.018900P PS=0.460000U PD=0.640000U
M_M2 N_Z_M7_d N_3_M7_g N_VSS_M6_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.018900P AD=0.033500P PS=0.640000U PD=0.830000U
M_M3 noxref_9 N_A_M8_g N_Z_M7_d VSS NMOS_VTL L=0.050U W=0.260000U AS=0.033500P AD=0.036400P PS=0.830000U PD=0.800000U
M_M4 N_VSS_M9_d N_B_M9_g noxref_9 VSS NMOS_VTL L=0.050U W=0.260000U AS=0.036400P AD=0.027300P PS=0.800000U PD=0.730000U
C_x_PM_XOR2_X2__VSS_c0 VSS x_PM_XOR2_X2__VSS_22 2.92244e-18
C_x_PM_XOR2_X2__VSS_c1 VSS N_VSS_M9_d 1.78745e-17
C_x_PM_XOR2_X2__VSS_c2 VSS x_PM_XOR2_X2__VSS_14 6.68756e-17
C_x_PM_XOR2_X2__VSS_c3 VSS N_VSS_M6_d 3.00222e-17
C_x_PM_XOR2_X2__VSS_c4 VSS x_PM_XOR2_X2__VSS_9 1.09715e-17
C_x_PM_XOR2_X2__VSS_c5 VSS x_PM_XOR2_X2__VSS_8 3.03506e-17
C_x_PM_XOR2_X2__VSS_c6 VSS N_VSS_M5_s 2.75676e-17
R_x_PM_XOR2_X2__VSS_r7 N_VSS_M9_d x_PM_XOR2_X2__VSS_18 0.230714
R_x_PM_XOR2_X2__VSS_r8 x_PM_XOR2_X2__VSS_22 x_PM_XOR2_X2__VSS_15 0.0731438
R_x_PM_XOR2_X2__VSS_r9 VSS x_PM_XOR2_X2__VSS_15 0.19
R_x_PM_XOR2_X2__VSS_r10 x_PM_XOR2_X2__VSS_18 x_PM_XOR2_X2__VSS_14 0.264221
R_x_PM_XOR2_X2__VSS_r11 VSS x_PM_XOR2_X2__VSS_14 0.961176
R_x_PM_XOR2_X2__VSS_r12 x_PM_XOR2_X2__VSS_22 x_PM_XOR2_X2__VSS_10 0.145286
R_x_PM_XOR2_X2__VSS_r13 N_VSS_M6_d x_PM_XOR2_X2__VSS_10 0.665
R_x_PM_XOR2_X2__VSS_r14 x_PM_XOR2_X2__VSS_22 x_PM_XOR2_X2__VSS_8 0.0731438
R_x_PM_XOR2_X2__VSS_r15 x_PM_XOR2_X2__VSS_9 x_PM_XOR2_X2__VSS_8 0.681765
R_x_PM_XOR2_X2__VSS_r16 x_PM_XOR2_X2__VSS_9 x_PM_XOR2_X2__VSS_4 0.264221
R_x_PM_XOR2_X2__VSS_r17 N_VSS_M5_s x_PM_XOR2_X2__VSS_4 0.665
C_x_PM_XOR2_X2__VDD_c0 VSS x_PM_XOR2_X2__VDD_11 5.06462e-17
C_x_PM_XOR2_X2__VDD_c1 VSS x_PM_XOR2_X2__VDD_8 9.04239e-17
C_x_PM_XOR2_X2__VDD_c2 VSS N_VDD_M1_d 1.60113e-17
R_x_PM_XOR2_X2__VDD_r3 x_PM_XOR2_X2__VDD_11 x_PM_XOR2_X2__VDD_8 0.0731438
R_x_PM_XOR2_X2__VDD_r4 VDD x_PM_XOR2_X2__VDD_8 0.178824
R_x_PM_XOR2_X2__VDD_r5 x_PM_XOR2_X2__VDD_11 x_PM_XOR2_X2__VDD_4 0.145286
R_x_PM_XOR2_X2__VDD_r6 N_VDD_M1_d x_PM_XOR2_X2__VDD_4 0.230714
C_x_PM_XOR2_X2__3_c0 VSS x_PM_XOR2_X2__3_32 1.23496e-17
C_x_PM_XOR2_X2__3_c1 VSS x_PM_XOR2_X2__3_24 2.62007e-17
C_x_PM_XOR2_X2__3_c2 VSS x_PM_XOR2_X2__3_23 5.632e-18
C_x_PM_XOR2_X2__3_c3 VSS x_PM_XOR2_X2__3_21 2.20346e-17
C_x_PM_XOR2_X2__3_c4 VSS N_3_M5_d 4.51028e-17
C_x_PM_XOR2_X2__3_c5 VSS x_PM_XOR2_X2__3_16 1.44792e-17
C_x_PM_XOR2_X2__3_c6 VSS x_PM_XOR2_X2__3_15 1.10108e-17
C_x_PM_XOR2_X2__3_c7 VSS N_3_M0_s 9.96232e-17
C_x_PM_XOR2_X2__3_c8 VSS N_3_M2_g 9.32321e-17
C_x_PM_XOR2_X2__3_c9 VSS N_3_M7_g 2.97214e-17
R_x_PM_XOR2_X2__3_r10 x_PM_XOR2_X2__3_32 x_PM_XOR2_X2__3_30 5.46
R_x_PM_XOR2_X2__3_r11 x_PM_XOR2_X2__3_30 x_PM_XOR2_X2__3_27 25.0012
R_x_PM_XOR2_X2__3_r12 x_PM_XOR2_X2__3_27 x_PM_XOR2_X2__3_24 0.176429
R_x_PM_XOR2_X2__3_r13 x_PM_XOR2_X2__3_23 x_PM_XOR2_X2__3_22 0.160909
R_x_PM_XOR2_X2__3_r14 x_PM_XOR2_X2__3_24 x_PM_XOR2_X2__3_21 0.095
R_x_PM_XOR2_X2__3_r15 x_PM_XOR2_X2__3_22 x_PM_XOR2_X2__3_21 0.895714
R_x_PM_XOR2_X2__3_r16 x_PM_XOR2_X2__3_23 x_PM_XOR2_X2__3_17 0.0418175
R_x_PM_XOR2_X2__3_r17 N_3_M5_d x_PM_XOR2_X2__3_17 0.800714
R_x_PM_XOR2_X2__3_r18 x_PM_XOR2_X2__3_23 x_PM_XOR2_X2__3_15 0.160909
R_x_PM_XOR2_X2__3_r19 x_PM_XOR2_X2__3_16 x_PM_XOR2_X2__3_15 0.624286
R_x_PM_XOR2_X2__3_r20 x_PM_XOR2_X2__3_16 x_PM_XOR2_X2__3_11 0.212645
R_x_PM_XOR2_X2__3_r21 N_3_M0_s x_PM_XOR2_X2__3_11 3.61
R_x_PM_XOR2_X2__3_r22 x_PM_XOR2_X2__3_32 x_PM_XOR2_X2__3_5 1.95
R_x_PM_XOR2_X2__3_r23 N_3_M2_g x_PM_XOR2_X2__3_5 99.84
R_x_PM_XOR2_X2__3_r24 x_PM_XOR2_X2__3_32 x_PM_XOR2_X2__3_VSS 1.95
R_x_PM_XOR2_X2__3_r25 N_3_M7_g x_PM_XOR2_X2__3_VSS 21.84
C_x_PM_XOR2_X2__A_c0 VSS x_PM_XOR2_X2__A_36 1.60834e-17
C_x_PM_XOR2_X2__A_c1 VSS x_PM_XOR2_X2__A_26 1.21081e-17
C_x_PM_XOR2_X2__A_c2 VSS x_PM_XOR2_X2__A_22 6.23618e-17
C_x_PM_XOR2_X2__A_c3 VSS x_PM_XOR2_X2__A_18 8.15108e-17
C_x_PM_XOR2_X2__A_c4 VSS N_A_M3_g 5.31977e-17
C_x_PM_XOR2_X2__A_c5 VSS N_A_M8_g 8.25873e-17
C_x_PM_XOR2_X2__A_c6 VSS N_A_M0_g 5.15027e-17
C_x_PM_XOR2_X2__A_c7 VSS N_A_M5_g 8.25861e-17
R_x_PM_XOR2_X2__A_r8 x_PM_XOR2_X2__A_26 x_PM_XOR2_X2__A_30 3.9
R_x_PM_XOR2_X2__A_r9 x_PM_XOR2_X2__A_26 x_PM_XOR2_X2__A_24 25.0012
R_x_PM_XOR2_X2__A_r10 A x_PM_XOR2_X2__A_24 0.124483
R_x_PM_XOR2_X2__A_r11 x_PM_XOR2_X2__A_24 x_PM_XOR2_X2__A_22 0.0851724
R_x_PM_XOR2_X2__A_r12 x_PM_XOR2_X2__A_36 x_PM_XOR2_X2__A_20 7.02
R_x_PM_XOR2_X2__A_r13 x_PM_XOR2_X2__A_20 x_PM_XOR2_X2__A_18 25.0012
R_x_PM_XOR2_X2__A_r14 x_PM_XOR2_X2__A_22 x_PM_XOR2_X2__A_17 0.095
R_x_PM_XOR2_X2__A_r15 x_PM_XOR2_X2__A_18 x_PM_XOR2_X2__A_17 1.995
R_x_PM_XOR2_X2__A_r16 x_PM_XOR2_X2__A_36 x_PM_XOR2_X2__A_13 1.95
R_x_PM_XOR2_X2__A_r17 N_A_M3_g x_PM_XOR2_X2__A_13 39
R_x_PM_XOR2_X2__A_r18 x_PM_XOR2_X2__A_36 x_PM_XOR2_X2__A_9 1.95
R_x_PM_XOR2_X2__A_r19 N_A_M8_g x_PM_XOR2_X2__A_9 88.92
R_x_PM_XOR2_X2__A_r20 x_PM_XOR2_X2__A_30 x_PM_XOR2_X2__A_5 1.95
R_x_PM_XOR2_X2__A_r21 N_A_M0_g x_PM_XOR2_X2__A_5 48.75
R_x_PM_XOR2_X2__A_r22 x_PM_XOR2_X2__A_30 x_PM_XOR2_X2__A_VSS 1.95
R_x_PM_XOR2_X2__A_r23 N_A_M5_g x_PM_XOR2_X2__A_VSS 95.16
C_x_PM_XOR2_X2__B_c0 VSS x_PM_XOR2_X2__B_35 1.25048e-17
C_x_PM_XOR2_X2__B_c1 VSS x_PM_XOR2_X2__B_24 8.22451e-18
C_x_PM_XOR2_X2__B_c2 VSS x_PM_XOR2_X2__B_22 3.95314e-17
C_x_PM_XOR2_X2__B_c3 VSS x_PM_XOR2_X2__B_18 1.2109e-16
C_x_PM_XOR2_X2__B_c4 VSS N_B_M4_g 6.79516e-17
C_x_PM_XOR2_X2__B_c5 VSS N_B_M9_g 6.48967e-17
C_x_PM_XOR2_X2__B_c6 VSS N_B_M1_g 7.2975e-17
C_x_PM_XOR2_X2__B_c7 VSS N_B_M6_g 5.17135e-17
R_x_PM_XOR2_X2__B_r8 x_PM_XOR2_X2__B_28 B 0.095
R_x_PM_XOR2_X2__B_r9 x_PM_XOR2_X2__B_32 x_PM_XOR2_X2__B_24 4.7687
R_x_PM_XOR2_X2__B_r10 x_PM_XOR2_X2__B_31 x_PM_XOR2_X2__B_24 4.7687
R_x_PM_XOR2_X2__B_r11 x_PM_XOR2_X2__B_24 x_PM_XOR2_X2__B_22 25.0012
R_x_PM_XOR2_X2__B_r12 B x_PM_XOR2_X2__B_22 0.00730769
R_x_PM_XOR2_X2__B_r13 x_PM_XOR2_X2__B_35 x_PM_XOR2_X2__B_20 4.42
R_x_PM_XOR2_X2__B_r14 x_PM_XOR2_X2__B_20 x_PM_XOR2_X2__B_18 25.0012
R_x_PM_XOR2_X2__B_r15 x_PM_XOR2_X2__B_28 x_PM_XOR2_X2__B_17 0.095
R_x_PM_XOR2_X2__B_r16 x_PM_XOR2_X2__B_18 x_PM_XOR2_X2__B_17 2.64733
R_x_PM_XOR2_X2__B_r17 x_PM_XOR2_X2__B_35 x_PM_XOR2_X2__B_13 1.95
R_x_PM_XOR2_X2__B_r18 N_B_M4_g x_PM_XOR2_X2__B_13 65.52
R_x_PM_XOR2_X2__B_r19 x_PM_XOR2_X2__B_35 x_PM_XOR2_X2__B_9 1.95
R_x_PM_XOR2_X2__B_r20 N_B_M9_g x_PM_XOR2_X2__B_9 62.4
R_x_PM_XOR2_X2__B_r21 N_B_M1_g x_PM_XOR2_X2__B_32 85.41
R_x_PM_XOR2_X2__B_r22 N_B_M6_g x_PM_XOR2_X2__B_31 58.5
C_x_PM_XOR2_X2__Z_c0 VSS x_PM_XOR2_X2__Z_16 2.93962e-17
C_x_PM_XOR2_X2__Z_c1 VSS x_PM_XOR2_X2__Z_14 2.66606e-17
C_x_PM_XOR2_X2__Z_c2 VSS x_PM_XOR2_X2__Z_13 2.89113e-17
C_x_PM_XOR2_X2__Z_c3 VSS Z 3.24504e-17
C_x_PM_XOR2_X2__Z_c4 VSS x_PM_XOR2_X2__Z_3 9.34374e-17
R_x_PM_XOR2_X2__Z_r5 x_PM_XOR2_X2__Z_16 x_PM_XOR2_X2__Z_15 1.87286
R_x_PM_XOR2_X2__Z_r6 x_PM_XOR2_X2__Z_16 x_PM_XOR2_X2__Z_13 0.212317
R_x_PM_XOR2_X2__Z_r7 x_PM_XOR2_X2__Z_14 x_PM_XOR2_X2__Z_13 0.787143
R_x_PM_XOR2_X2__Z_r8 N_Z_M3_d Z 0.257857
R_x_PM_XOR2_X2__Z_r9 x_PM_XOR2_X2__Z_14 x_PM_XOR2_X2__Z_7 0.212317
R_x_PM_XOR2_X2__Z_r10 Z x_PM_XOR2_X2__Z_7 0.407143
R_x_PM_XOR2_X2__Z_r11 x_PM_XOR2_X2__Z_15 x_PM_XOR2_X2__Z_3 0.244544
R_x_PM_XOR2_X2__Z_r12 N_Z_M7_d x_PM_XOR2_X2__Z_3 1.01107
C_x_PM_XOR2_X2__7_c0 VSS N_7_M4_d 7.56582e-17
R_x_PM_XOR2_X2__7_r1 N_7_M4_d N_7_M2_d 2.03571
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
