.SUBCKT or2 A1 A2 VDD VSS ZN 
M_M3 7 N_A1_M0_g N_3_M0_s VDD PMOS_VTL L=0.050U W=0.195000U AS=0.020475P AD=0.027300P PS=0.600000U PD=0.670000U
M_M4 N_VDD_M1_d N_A2_M1_g 7 VDD PMOS_VTL L=0.050U W=0.195000U AS=0.027300P AD=0.037950P PS=0.670000U PD=0.860000U
M_M5 N_ZN_M2_d N_3_M2_g N_VDD_M1_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037950P AD=0.028350P PS=0.860000U PD=0.750000U
M_M0 N_3_M3_d N_A1_M3_g N_VSS_M3_s VSS NMOS_VTL L=0.050U W=0.090000U AS=0.009450P AD=0.012600P PS=0.390000U PD=0.460000U
M_M1 N_VSS_M4_d N_A2_M4_g N_3_M3_d VSS NMOS_VTL L=0.050U W=0.090000U AS=0.012600P AD=0.023850P PS=0.460000U PD=0.680000U
M_M2 N_ZN_M5_d N_3_M5_g N_VSS_M4_d VSS NMOS_VTL L=0.050U W=0.180000U AS=0.023850P AD=0.018900P PS=0.680000U PD=0.570000U
C_x_PM_OR2_X2__VSS_c0 VSS x_PM_OR2_X2__VSS_15 3.72032e-17
C_x_PM_OR2_X2__VSS_c1 VSS N_VSS_M4_d 1.48795e-17
C_x_PM_OR2_X2__VSS_c2 VSS x_PM_OR2_X2__VSS_6 1.07612e-17
C_x_PM_OR2_X2__VSS_c3 VSS x_PM_OR2_X2__VSS_5 3.45483e-17
C_x_PM_OR2_X2__VSS_c4 VSS x_PM_OR2_X2__VSS_4 2.26908e-17
R_x_PM_OR2_X2__VSS_r5 x_PM_OR2_X2__VSS_15 x_PM_OR2_X2__VSS_9 0.145286
R_x_PM_OR2_X2__VSS_r6 N_VSS_M4_d x_PM_OR2_X2__VSS_9 0.230714
R_x_PM_OR2_X2__VSS_r7 VSS x_PM_OR2_X2__VSS_6 0.603529
R_x_PM_OR2_X2__VSS_r8 x_PM_OR2_X2__VSS_15 x_PM_OR2_X2__VSS_5 0.0731438
R_x_PM_OR2_X2__VSS_r9 VSS x_PM_OR2_X2__VSS_5 0.134118
R_x_PM_OR2_X2__VSS_r10 x_PM_OR2_X2__VSS_6 x_PM_OR2_X2__VSS_4 0.264221
R_x_PM_OR2_X2__VSS_r11 x_PM_OR2_X2__VSS_4 N_VSS_M3_s 0.543196
C_x_PM_OR2_X2__VDD_c0 VSS x_PM_OR2_X2__VDD_12 4.05231e-17
C_x_PM_OR2_X2__VDD_c1 VSS N_VDD_M1_d 2.06356e-17
C_x_PM_OR2_X2__VDD_c2 VSS x_PM_OR2_X2__VDD_2 4.07936e-17
R_x_PM_OR2_X2__VDD_r3 x_PM_OR2_X2__VDD_12 x_PM_OR2_X2__VDD_6 0.145286
R_x_PM_OR2_X2__VDD_r4 N_VDD_M1_d x_PM_OR2_X2__VDD_6 0.420714
R_x_PM_OR2_X2__VDD_r5 x_PM_OR2_X2__VDD_12 x_PM_OR2_X2__VDD_2 0.0731438
R_x_PM_OR2_X2__VDD_r6 VDD x_PM_OR2_X2__VDD_2 0.0782353
C_x_PM_OR2_X2__3_c0 VSS x_PM_OR2_X2__3_31 1.75553e-17
C_x_PM_OR2_X2__3_c1 VSS x_PM_OR2_X2__3_28 1.72947e-17
C_x_PM_OR2_X2__3_c2 VSS x_PM_OR2_X2__3_25 5.24935e-17
C_x_PM_OR2_X2__3_c3 VSS x_PM_OR2_X2__3_22 2.8529e-17
C_x_PM_OR2_X2__3_c4 VSS N_3_M3_d 4.52149e-17
C_x_PM_OR2_X2__3_c5 VSS x_PM_OR2_X2__3_16 1.69957e-17
C_x_PM_OR2_X2__3_c6 VSS x_PM_OR2_X2__3_15 3.68802e-17
C_x_PM_OR2_X2__3_c7 VSS N_3_M0_s 4.3344e-17
C_x_PM_OR2_X2__3_c8 VSS N_3_M2_g 9.38216e-17
C_x_PM_OR2_X2__3_c9 VSS N_3_M5_g 4.44376e-17
R_x_PM_OR2_X2__3_r10 x_PM_OR2_X2__3_31 x_PM_OR2_X2__3_29 7.54
R_x_PM_OR2_X2__3_r11 x_PM_OR2_X2__3_29 x_PM_OR2_X2__3_25 25.0012
R_x_PM_OR2_X2__3_r12 x_PM_OR2_X2__3_28 x_PM_OR2_X2__3_23 0.0418175
R_x_PM_OR2_X2__3_r13 x_PM_OR2_X2__3_25 x_PM_OR2_X2__3_23 1.045
R_x_PM_OR2_X2__3_r14 x_PM_OR2_X2__3_28 x_PM_OR2_X2__3_21 0.160909
R_x_PM_OR2_X2__3_r15 x_PM_OR2_X2__3_22 x_PM_OR2_X2__3_21 0.705714
R_x_PM_OR2_X2__3_r16 x_PM_OR2_X2__3_28 x_PM_OR2_X2__3_17 0.160909
R_x_PM_OR2_X2__3_r17 N_3_M3_d x_PM_OR2_X2__3_17 1.045
R_x_PM_OR2_X2__3_r18 x_PM_OR2_X2__3_22 x_PM_OR2_X2__3_15 0.212317
R_x_PM_OR2_X2__3_r19 x_PM_OR2_X2__3_16 x_PM_OR2_X2__3_15 0.651429
R_x_PM_OR2_X2__3_r20 x_PM_OR2_X2__3_16 x_PM_OR2_X2__3_11 0.212317
R_x_PM_OR2_X2__3_r21 N_3_M0_s x_PM_OR2_X2__3_11 2.29357
R_x_PM_OR2_X2__3_r22 x_PM_OR2_X2__3_31 x_PM_OR2_X2__3_5 1.95
R_x_PM_OR2_X2__3_r23 N_3_M2_g x_PM_OR2_X2__3_5 99.84
R_x_PM_OR2_X2__3_r24 x_PM_OR2_X2__3_31 x_PM_OR2_X2__3_VSS 1.95
R_x_PM_OR2_X2__3_r25 N_3_M5_g x_PM_OR2_X2__3_VSS 38.22
C_x_PM_OR2_X2__A1_c0 VSS x_PM_OR2_X2__A1_18 8.81315e-18
C_x_PM_OR2_X2__A1_c1 VSS x_PM_OR2_X2__A1_12 5.4822e-17
C_x_PM_OR2_X2__A1_c2 VSS N_A1_M0_g 8.90209e-17
C_x_PM_OR2_X2__A1_c3 VSS N_A1_M3_g 3.57915e-17
R_x_PM_OR2_X2__A1_r4 x_PM_OR2_X2__A1_18 x_PM_OR2_X2__A1_14 3.38
R_x_PM_OR2_X2__A1_r5 x_PM_OR2_X2__A1_14 x_PM_OR2_X2__A1_12 25.0012
R_x_PM_OR2_X2__A1_r6 x_PM_OR2_X2__A1_12 A1 0.115357
R_x_PM_OR2_X2__A1_r7 x_PM_OR2_X2__A1_18 x_PM_OR2_X2__A1_5 1.95
R_x_PM_OR2_X2__A1_r8 N_A1_M0_g x_PM_OR2_X2__A1_5 101.01
R_x_PM_OR2_X2__A1_r9 x_PM_OR2_X2__A1_18 x_PM_OR2_X2__A1_VSS 1.95
R_x_PM_OR2_X2__A1_r10 N_A1_M3_g x_PM_OR2_X2__A1_VSS 35.88
C_x_PM_OR2_X2__A2_c0 VSS A2 6.95827e-17
C_x_PM_OR2_X2__A2_c1 VSS x_PM_OR2_X2__A2_11 1.12977e-17
C_x_PM_OR2_X2__A2_c2 VSS N_A2_M1_g 6.44459e-17
C_x_PM_OR2_X2__A2_c3 VSS N_A2_M4_g 5.20861e-17
R_x_PM_OR2_X2__A2_r4 x_PM_OR2_X2__A2_11 x_PM_OR2_X2__A2_16 4.42
R_x_PM_OR2_X2__A2_r5 x_PM_OR2_X2__A2_11 x_PM_OR2_X2__A2_9 25.0012
R_x_PM_OR2_X2__A2_r6 A2 x_PM_OR2_X2__A2_9 0.196786
R_x_PM_OR2_X2__A2_r7 x_PM_OR2_X2__A2_16 x_PM_OR2_X2__A2_5 1.95
R_x_PM_OR2_X2__A2_r8 N_A2_M1_g x_PM_OR2_X2__A2_5 79.95
R_x_PM_OR2_X2__A2_r9 x_PM_OR2_X2__A2_16 x_PM_OR2_X2__A2_VSS 1.95
R_x_PM_OR2_X2__A2_r10 N_A2_M4_g x_PM_OR2_X2__A2_VSS 56.94
C_x_PM_OR2_X2__ZN_c0 VSS N_ZN_M5_d 1.3351e-16
R_x_PM_OR2_X2__ZN_r1 N_ZN_M2_d ZN 2.23929
R_x_PM_OR2_X2__ZN_r2 ZN N_ZN_M5_d 2.91786
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
