.SUBCKT oai3 B1 B2 A VDD VSS ZN 
M_M3 noxref_8 N_B2_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.390000U AS=0.040950P AD=0.054600P PS=0.990000U PD=1.060000U
M_M4 N_ZN_M1_d N_B1_M1_g noxref_8 VDD PMOS_VTL L=0.050U W=0.390000U AS=0.054600P AD=0.046200P PS=1.060000U PD=1.060000U
M_M5 N_VDD_M2_d N_A_M2_g N_ZN_M1_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.046200P AD=0.028350P PS=1.060000U PD=0.750000U
M_M0 N_ZN_M3_d N_B2_M3_g N_3_M3_s VSS NMOS_VTL L=0.050U W=0.260000U AS=0.027300P AD=0.036400P PS=0.730000U PD=0.800000U
M_M1 N_3_M4_d N_B1_M4_g N_ZN_M3_d VSS NMOS_VTL L=0.050U W=0.260000U AS=0.036400P AD=0.036400P PS=0.800000U PD=0.800000U
M_M2 N_VSS_M5_d N_A_M5_g N_3_M4_d VSS NMOS_VTL L=0.050U W=0.260000U AS=0.036400P AD=0.027300P PS=0.800000U PD=0.730000U
C_x_PM_OAI21_X2__VSS_c0 VSS N_VSS_M5_d 2.20348e-17
C_x_PM_OAI21_X2__VSS_c1 VSS x_PM_OAI21_X2__VSS_2 1.54775e-16
R_x_PM_OAI21_X2__VSS_r2 N_VSS_M5_d x_PM_OAI21_X2__VSS_6 0.447857
R_x_PM_OAI21_X2__VSS_r3 x_PM_OAI21_X2__VSS_6 x_PM_OAI21_X2__VSS_2 0.264221
R_x_PM_OAI21_X2__VSS_r4 VSS x_PM_OAI21_X2__VSS_2 0.558824
C_x_PM_OAI21_X2__VDD_c0 VSS VDD 1.24485e-17
C_x_PM_OAI21_X2__VDD_c1 VSS N_VDD_M2_d 3.14319e-17
C_x_PM_OAI21_X2__VDD_c2 VSS x_PM_OAI21_X2__VDD_7 6.1596e-17
C_x_PM_OAI21_X2__VDD_c3 VSS N_VDD_M0_s 2.3501e-17
R_x_PM_OAI21_X2__VDD_r4 x_PM_OAI21_X2__VDD_16 VDD 0.225185
R_x_PM_OAI21_X2__VDD_r5 x_PM_OAI21_X2__VDD_15 VDD 0.101823
R_x_PM_OAI21_X2__VDD_r6 N_VDD_M2_d x_PM_OAI21_X2__VDD_9 0.420714
R_x_PM_OAI21_X2__VDD_r7 x_PM_OAI21_X2__VDD_16 x_PM_OAI21_X2__VDD_8 0.095
R_x_PM_OAI21_X2__VDD_r8 x_PM_OAI21_X2__VDD_9 x_PM_OAI21_X2__VDD_7 0.264221
R_x_PM_OAI21_X2__VDD_r9 x_PM_OAI21_X2__VDD_8 x_PM_OAI21_X2__VDD_7 1.10647
R_x_PM_OAI21_X2__VDD_r10 N_VDD_M0_s x_PM_OAI21_X2__VDD_15 0.420714
C_x_PM_OAI21_X2__3_c0 VSS N_3_M4_d 1.36966e-16
R_x_PM_OAI21_X2__3_r1 N_3_M4_d N_3_M3_s 2.03571
C_x_PM_OAI21_X2__B2_c0 VSS x_PM_OAI21_X2__B2_18 8.8921e-18
C_x_PM_OAI21_X2__B2_c1 VSS x_PM_OAI21_X2__B2_12 3.8522e-17
C_x_PM_OAI21_X2__B2_c2 VSS N_B2_M0_g 7.84586e-17
C_x_PM_OAI21_X2__B2_c3 VSS N_B2_M3_g 3.85693e-17
R_x_PM_OAI21_X2__B2_r4 x_PM_OAI21_X2__B2_18 x_PM_OAI21_X2__B2_14 4.42
R_x_PM_OAI21_X2__B2_r5 x_PM_OAI21_X2__B2_14 x_PM_OAI21_X2__B2_12 25.0012
R_x_PM_OAI21_X2__B2_r6 x_PM_OAI21_X2__B2_12 B2 0.156071
R_x_PM_OAI21_X2__B2_r7 x_PM_OAI21_X2__B2_18 x_PM_OAI21_X2__B2_5 1.95
R_x_PM_OAI21_X2__B2_r8 N_B2_M0_g x_PM_OAI21_X2__B2_5 85.8
R_x_PM_OAI21_X2__B2_r9 x_PM_OAI21_X2__B2_18 x_PM_OAI21_X2__B2_VSS 1.95
R_x_PM_OAI21_X2__B2_r10 N_B2_M3_g x_PM_OAI21_X2__B2_VSS 30.42
C_x_PM_OAI21_X2__ZN_c0 VSS N_ZN_M1_d 4.25468e-17
C_x_PM_OAI21_X2__ZN_c1 VSS x_PM_OAI21_X2__ZN_10 9.63135e-18
C_x_PM_OAI21_X2__ZN_c2 VSS x_PM_OAI21_X2__ZN_9 1.9166e-17
C_x_PM_OAI21_X2__ZN_c3 VSS N_ZN_M3_d 1.33496e-16
R_x_PM_OAI21_X2__ZN_r4 N_ZN_M1_d x_PM_OAI21_X2__ZN_11 0.746429
R_x_PM_OAI21_X2__ZN_r5 x_PM_OAI21_X2__ZN_11 x_PM_OAI21_X2__ZN_9 0.212317
R_x_PM_OAI21_X2__ZN_r6 x_PM_OAI21_X2__ZN_10 x_PM_OAI21_X2__ZN_9 0.651429
R_x_PM_OAI21_X2__ZN_r7 ZN N_ZN_M3_d 3.02643
R_x_PM_OAI21_X2__ZN_r8 x_PM_OAI21_X2__ZN_10 x_PM_OAI21_X2__ZN_3 0.212317
R_x_PM_OAI21_X2__ZN_r9 ZN x_PM_OAI21_X2__ZN_3 0.352857
C_x_PM_OAI21_X2__B1_c0 VSS B1 6.15349e-17
C_x_PM_OAI21_X2__B1_c1 VSS x_PM_OAI21_X2__B1_11 1.04443e-17
C_x_PM_OAI21_X2__B1_c2 VSS N_B1_M1_g 8.33914e-17
C_x_PM_OAI21_X2__B1_c3 VSS N_B1_M4_g 4.15528e-17
R_x_PM_OAI21_X2__B1_r4 x_PM_OAI21_X2__B1_11 x_PM_OAI21_X2__B1_16 3.38
R_x_PM_OAI21_X2__B1_r5 x_PM_OAI21_X2__B1_11 x_PM_OAI21_X2__B1_9 25.0012
R_x_PM_OAI21_X2__B1_r6 B1 x_PM_OAI21_X2__B1_9 0.156071
R_x_PM_OAI21_X2__B1_r7 x_PM_OAI21_X2__B1_16 x_PM_OAI21_X2__B1_5 1.95
R_x_PM_OAI21_X2__B1_r8 N_B1_M1_g x_PM_OAI21_X2__B1_5 86.58
R_x_PM_OAI21_X2__B1_r9 x_PM_OAI21_X2__B1_16 x_PM_OAI21_X2__B1_VSS 1.95
R_x_PM_OAI21_X2__B1_r10 N_B1_M4_g x_PM_OAI21_X2__B1_VSS 29.64
C_x_PM_OAI21_X2__A_c0 VSS A 3.72975e-17
C_x_PM_OAI21_X2__A_c1 VSS x_PM_OAI21_X2__A_11 8.36959e-18
C_x_PM_OAI21_X2__A_c2 VSS N_A_M2_g 7.78115e-17
C_x_PM_OAI21_X2__A_c3 VSS N_A_M5_g 3.90983e-17
R_x_PM_OAI21_X2__A_r4 x_PM_OAI21_X2__A_11 x_PM_OAI21_X2__A_16 3.38
R_x_PM_OAI21_X2__A_r5 x_PM_OAI21_X2__A_11 x_PM_OAI21_X2__A_9 25.0012
R_x_PM_OAI21_X2__A_r6 A x_PM_OAI21_X2__A_9 0.156071
R_x_PM_OAI21_X2__A_r7 x_PM_OAI21_X2__A_16 x_PM_OAI21_X2__A_5 1.95
R_x_PM_OAI21_X2__A_r8 N_A_M2_g x_PM_OAI21_X2__A_5 95.16
R_x_PM_OAI21_X2__A_r9 x_PM_OAI21_X2__A_16 x_PM_OAI21_X2__A_VSS 1.95
R_x_PM_OAI21_X2__A_r10 N_A_M5_g x_PM_OAI21_X2__A_VSS 30.42
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
