module singlepath (N4, N2892);
input N4;
output N2892;
wire N2873, N2846, N2828, N2810, N2809, N2776, N2750, N1999, N1958, N1310, N1879, N346, N1774, N2000, N1849, N1823, N1709, N1708, N1651, N2651, N1824, N2573, N559, N1443, N2606, N1944, N2078, N1208, N1647, N1010, N2648, N2874, N1013, N2020, N1207, N1513, N634, N2642, N194, N1546, N1487, N1444, N2038, N2060, N2196, N1355, N2199, N2224, N2627, N2570, N2225, N2297, N2549, N2645, N2233, N1746, N2241, N2263, N2266, N2552, N2286, N2555, N2576, N2597, N2600, N2603, N2746, Vcc, gnd;
not NOT1_2(N194, N4);
buf BUFF1_44(N346, N4);
buf BUFF1_82(N559, N194);
buf BUFF1_107(N634, N194);
buf BUFF1_219(N1010, N559);
buf BUFF1_220(N1013, N559);
not NOT1_272(N1207, N1013);
nand NAND2_273(N1208, N1013, Vcc);
nand NAND2_314(N1310, N1207, Vcc);
nand NAND2_336(N1355, N1310, Vcc);
nand NAND2_366(N1443, N1355, Vcc);
not NOT1_367(N1444, N1355);
nand NAND2_396(N1487, N1444, Vcc);
nand NAND2_412(N1513, N1487, Vcc);
not NOT1_428(N1546, N1513);
buf BUFF1_457(N1647, N1546);
buf BUFF1_458(N1651, N1546);
nand NAND2_478(N1708, N1647, Vcc);
not NOT1_479(N1709, N1647);
nand NAND2_497(N1746, N1709, Vcc);
nand NAND2_510(N1774, N1746, Vcc);
nand NAND2_534(N1823, N1774, Vcc);
not NOT1_535(N1824, N1774);
nand NAND2_544(N1849, N1824, Vcc);
nand NAND2_558(N1879, N1849, Vcc);
buf BUFF1_588(N1944, N1879);
buf BUFF1_592(N1958, N1879);
not NOT1_604(N1999, N1944);
nand NAND2_605(N2000, N1944, Vcc);
nand NAND2_621(N2020, N1999, Vcc);
nand NAND2_633(N2038, N2020, Vcc);
not NOT1_641(N2060, N2038);
nand NAND2_649(N2078, N2060, Vcc);
buf BUFF1_659(N2196, N2078);
buf BUFF1_660(N2199, N2078);
nand NAND2_669(N2224, N2196, Vcc);
not NOT1_670(N2225, N2196);
nand NAND2_678(N2233, N2225, Vcc);
nand NAND2_684(N2241, N2233, Vcc);
not NOT1_692(N2263, N2241);
and AND2_693(N2266, N2241, Vcc);
buf BUFF1_697(N2286, N2266);
buf BUFF1_698(N2297, N2266);
nand NAND5_714(N2549, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_715(N2552, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_716(N2555, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_721(N2570, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_722(N2573, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_723(N2576, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_725(N2597, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_726(N2600, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_727(N2603, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_728(N2606, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND5_733(N2627, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_742(N2642, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_743(N2645, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_744(N2648, N2297, Vcc, Vcc, Vcc, Vcc);
and AND5_745(N2651, N2297, Vcc, Vcc, Vcc, Vcc);
nand NAND8_791(N2746, N2555, Vcc, Vcc, Vcc, Vcc, Vcc, Vcc, Vcc);
and AND8_793(N2750, N2555, Vcc, Vcc, Vcc, Vcc, Vcc, Vcc, Vcc);
and AND2_811(N2776, N2746, Vcc);
nand NAND2_826(N2809, N2776, Vcc);
not NOT1_827(N2810, N2776);
nand NAND2_835(N2828, N2810, Vcc);
nand NAND2_838(N2846, N2828, Vcc);
nand NAND2_858(N2873, N2846, Vcc);
not NOT1_859(N2874, N2846);
nand NAND2_875(N2892, N2873, Vcc);

endmodule
