.SUBCKT nand2 A1 A2 VDD VSS ZN 
M_M2 N_ZN_M0_d N_A2_M0_g N_VDD_M0_s VDD PMOS_VTL L=0.050U W=0.270000U AS=0.028350P AD=0.037800P PS=0.750000U PD=0.820000U
M_M3 N_VDD_M1_d N_A1_M1_g N_ZN_M0_d VDD PMOS_VTL L=0.050U W=0.270000U AS=0.037800P AD=0.028350P PS=0.820000U PD=0.750000U
M_M0 6 N_A2_M2_g N_VSS_M2_s VSS NMOS_VTL L=0.050U W=0.260000U AS=0.027300P AD=0.036400P PS=0.730000U PD=0.800000U
M_M1 N_ZN_M3_d N_A1_M3_g 6 VSS NMOS_VTL L=0.050U W=0.260000U AS=0.036400P AD=0.027300P PS=0.800000U PD=0.730000U
C_x_PM_NAND2_X2__VSS_c0 VSS VSS 5.03826e-17
C_x_PM_NAND2_X2__VSS_c1 VSS x_PM_NAND2_X2__VSS_6 1.04465e-17
C_x_PM_NAND2_X2__VSS_c2 VSS N_VSS_M2_s 1.83058e-17
R_x_PM_NAND2_X2__VSS_r3 VSS x_PM_NAND2_X2__VSS_6 0.391176
R_x_PM_NAND2_X2__VSS_r4 x_PM_NAND2_X2__VSS_6 x_PM_NAND2_X2__VSS_2 0.264221
R_x_PM_NAND2_X2__VSS_r5 N_VSS_M2_s x_PM_NAND2_X2__VSS_2 0.230714
C_x_PM_NAND2_X2__VDD_c0 VSS N_VDD_M1_d 4.75732e-17
C_x_PM_NAND2_X2__VDD_c1 VSS x_PM_NAND2_X2__VDD_7 4.67275e-17
C_x_PM_NAND2_X2__VDD_c2 VSS N_VDD_M0_s 2.99432e-17
C_x_PM_NAND2_X2__VDD_c3 VSS x_PM_NAND2_X2__VDD_3 1.06496e-17
R_x_PM_NAND2_X2__VDD_r4 N_VDD_M1_d x_PM_NAND2_X2__VDD_9 0.420714
R_x_PM_NAND2_X2__VDD_r5 VDD x_PM_NAND2_X2__VDD_8 0.195294
R_x_PM_NAND2_X2__VDD_r6 x_PM_NAND2_X2__VDD_9 x_PM_NAND2_X2__VDD_7 0.264221
R_x_PM_NAND2_X2__VDD_r7 x_PM_NAND2_X2__VDD_8 x_PM_NAND2_X2__VDD_7 0.681765
R_x_PM_NAND2_X2__VDD_r8 VDD x_PM_NAND2_X2__VDD_3 0.0689273
R_x_PM_NAND2_X2__VDD_r9 N_VDD_M0_s x_PM_NAND2_X2__VDD_3 0.420714
C_x_PM_NAND2_X2__A2_c0 VSS x_PM_NAND2_X2__A2_14 7.51478e-18
C_x_PM_NAND2_X2__A2_c1 VSS A2 6.01437e-17
C_x_PM_NAND2_X2__A2_c2 VSS N_A2_M0_g 8.26414e-17
C_x_PM_NAND2_X2__A2_c3 VSS N_A2_M2_g 3.58741e-17
R_x_PM_NAND2_X2__A2_r4 x_PM_NAND2_X2__A2_18 x_PM_NAND2_X2__A2_14 4.74714
R_x_PM_NAND2_X2__A2_r5 x_PM_NAND2_X2__A2_17 x_PM_NAND2_X2__A2_14 4.74714
R_x_PM_NAND2_X2__A2_r6 x_PM_NAND2_X2__A2_14 x_PM_NAND2_X2__A2_12 25.0012
R_x_PM_NAND2_X2__A2_r7 x_PM_NAND2_X2__A2_12 A2 0.266
R_x_PM_NAND2_X2__A2_r8 N_A2_M0_g x_PM_NAND2_X2__A2_18 103.74
R_x_PM_NAND2_X2__A2_r9 N_A2_M2_g x_PM_NAND2_X2__A2_17 28.08
C_x_PM_NAND2_X2__ZN_c0 VSS N_ZN_M3_d 9.46701e-17
C_x_PM_NAND2_X2__ZN_c1 VSS x_PM_NAND2_X2__ZN_8 7.68686e-18
C_x_PM_NAND2_X2__ZN_c2 VSS x_PM_NAND2_X2__ZN_7 3.24105e-17
C_x_PM_NAND2_X2__ZN_c3 VSS N_ZN_M0_d 6.2878e-17
R_x_PM_NAND2_X2__ZN_r4 ZN N_ZN_M3_d 1.93167
R_x_PM_NAND2_X2__ZN_r5 ZN x_PM_NAND2_X2__ZN_9 0.527778
R_x_PM_NAND2_X2__ZN_r6 x_PM_NAND2_X2__ZN_9 x_PM_NAND2_X2__ZN_7 0.21666
R_x_PM_NAND2_X2__ZN_r7 x_PM_NAND2_X2__ZN_8 x_PM_NAND2_X2__ZN_7 0.624286
R_x_PM_NAND2_X2__ZN_r8 x_PM_NAND2_X2__ZN_8 x_PM_NAND2_X2__ZN_3 0.212317
R_x_PM_NAND2_X2__ZN_r9 N_ZN_M0_d x_PM_NAND2_X2__ZN_3 1.18071
C_x_PM_NAND2_X2__A1_c0 VSS x_PM_NAND2_X2__A1_18 1.23667e-17
C_x_PM_NAND2_X2__A1_c1 VSS A1 8.87208e-17
C_x_PM_NAND2_X2__A1_c2 VSS N_A1_M1_g 9.96411e-17
C_x_PM_NAND2_X2__A1_c3 VSS N_A1_M3_g 3.7962e-17
R_x_PM_NAND2_X2__A1_r4 x_PM_NAND2_X2__A1_18 x_PM_NAND2_X2__A1_14 3.9
R_x_PM_NAND2_X2__A1_r5 x_PM_NAND2_X2__A1_14 x_PM_NAND2_X2__A1_12 25.0012
R_x_PM_NAND2_X2__A1_r6 x_PM_NAND2_X2__A1_12 A1 0.316667
R_x_PM_NAND2_X2__A1_r7 x_PM_NAND2_X2__A1_18 x_PM_NAND2_X2__A1_5 1.95
R_x_PM_NAND2_X2__A1_r8 N_A1_M1_g x_PM_NAND2_X2__A1_5 103.74
R_x_PM_NAND2_X2__A1_r9 x_PM_NAND2_X2__A1_18 x_PM_NAND2_X2__A1_VSS 1.95
R_x_PM_NAND2_X2__A1_r10 N_A1_M3_g x_PM_NAND2_X2__A1_VSS 28.08
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
